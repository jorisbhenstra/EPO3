configuration d_ff_behaviour_cfg of d_ff is
   for behaviour
   end for;
end d_ff_behaviour_cfg;
