configuration y_decider_behaviour_cfg of y_decider is
   for behaviour
   end for;
end y_decider_behaviour_cfg;
