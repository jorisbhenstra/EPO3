
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture synthesised of gradius_toplvl is

  component movement
    port(clk           : in  std_logic;
         reset         : in  std_logic;
         frame_ready   : in  std_logic;
         left          : in  std_logic;
         right         : in  std_logic;
         up            : in  std_logic;
         down          : in  std_logic;
         shoot         : in  std_logic;
         enemy_1_y     : in  std_logic_vector(8 downto 0);
         enemy_2_y     : in  std_logic_vector(8 downto 0);
         enemy_3_y     : in  std_logic_vector(8 downto 0);
         enemy_4_y     : in  std_logic_vector(8 downto 0);
         enemy_5_y     : in  std_logic_vector(8 downto 0);
         enemy_6_y     : in  std_logic_vector(8 downto 0);
         e_respawn_1   : in  std_logic;
         e_respawn_2   : in  std_logic;
         e_respawn_3   : in  std_logic;
         e_respawn_4   : in  std_logic;
         e_respawn_5   : in  std_logic;
         e_respawn_6   : in  std_logic;
         coll_enemy_1  : in  std_logic;
         coll_enemy_2  : in  std_logic;
         coll_enemy_3  : in  std_logic;
         coll_enemy_4  : in  std_logic;
         coll_enemy_5  : in  std_logic;
         coll_enemy_6  : in  std_logic;
         coll_bullet_1 : in  std_logic;
         coll_bullet_2 : in  std_logic;
         coll_bullet_3 : in  std_logic;
         coll_player   : in  std_logic;
         player_x      : out std_logic_vector(8 downto 0);
         player_y      : out std_logic_vector(8 downto 0);
         enemy_x_1     : out std_logic_vector(8 downto 0);
         enemy_y_1     : out std_logic_vector(8 downto 0);
         enemy_x_2     : out std_logic_vector(8 downto 0);
         enemy_y_2     : out std_logic_vector(8 downto 0);
         enemy_x_3     : out std_logic_vector(8 downto 0);
         enemy_y_3     : out std_logic_vector(8 downto 0);
         enemy_x_4     : out std_logic_vector(8 downto 0);
         enemy_y_4     : out std_logic_vector(8 downto 0);
         enemy_x_5     : out std_logic_vector(8 downto 0);
         enemy_y_5     : out std_logic_vector(8 downto 0);
         enemy_x_6     : out std_logic_vector(8 downto 0);
         enemy_y_6     : out std_logic_vector(8 downto 0);
         bullet_x_1    : out std_logic_vector(8 downto 0);
         bullet_y_1    : out std_logic_vector(8 downto 0);
         bullet_x_2    : out std_logic_vector(8 downto 0);
         bullet_y_2    : out std_logic_vector(8 downto 0);
         bullet_x_3    : out std_logic_vector(8 downto 0);
         bullet_y_3    : out std_logic_vector(8 downto 0);
         enemy_alive_1 : out std_logic;
         enemy_alive_2 : out std_logic;
         enemy_alive_3 : out std_logic;
         enemy_alive_4 : out std_logic;
         enemy_alive_5 : out std_logic;
         enemy_alive_6 : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component ND2D4BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component AO31D0BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component AOI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AO32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IINR4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component MAOI222D0BWP7T
    port(A, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OA221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component AO222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component MUX2ND0BWP7T
    port(I0, I1, S : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component DFKSND1BWP7T
    port(CP, D, SN : in std_logic; Q, QN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component DFXQD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component DFCNQD1BWP7T
    port(CDN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component OAI33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OR3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component XNR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component OA32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component CKXOR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OA31D0BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component DFND1BWP7T
    port(CPN, D : in std_logic; Q, QN : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component HA1D0BWP7T
    port(A, B : in std_logic; CO, S : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CP, CN, D : in std_logic; Q, QN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component IOA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CP, CN, D : in std_logic; Q : out std_logic);
  end component;

  signal y_e_spawn_1 : std_logic_vector(8 downto 0);
  signal y_e_spawn_2 : std_logic_vector(8 downto 0);
  signal y_e_spawn_3 : std_logic_vector(8 downto 0);
  signal y_e_spawn_4 : std_logic_vector(8 downto 0);
  signal y_e_spawn_5 : std_logic_vector(8 downto 0);
  signal collision_output_vector : std_logic_vector(15 downto 0);
  signal x_pos_p : std_logic_vector(8 downto 0);
  signal y_pos_p : std_logic_vector(8 downto 0);
  signal x_pos_e1 : std_logic_vector(8 downto 0);
  signal y_pos_e1 : std_logic_vector(8 downto 0);
  signal x_pos_e2 : std_logic_vector(8 downto 0);
  signal y_pos_e2 : std_logic_vector(8 downto 0);
  signal x_pos_e3 : std_logic_vector(8 downto 0);
  signal y_pos_e3 : std_logic_vector(8 downto 0);
  signal x_pos_e4 : std_logic_vector(8 downto 0);
  signal y_pos_e4 : std_logic_vector(8 downto 0);
  signal x_pos_e5 : std_logic_vector(8 downto 0);
  signal y_pos_e5 : std_logic_vector(8 downto 0);
  signal x_pos_e6 : std_logic_vector(8 downto 0);
  signal y_pos_e6 : std_logic_vector(8 downto 0);
  signal x_pos_b1 : std_logic_vector(8 downto 0);
  signal y_pos_b1 : std_logic_vector(8 downto 0);
  signal x_pos_b2 : std_logic_vector(8 downto 0);
  signal y_pos_b2 : std_logic_vector(8 downto 0);
  signal x_pos_b3 : std_logic_vector(8 downto 0);
  signal y_pos_b3 : std_logic_vector(8 downto 0);
  signal VGA_y : std_logic_vector(9 downto 0);
  signal VGA_x : std_logic_vector(8 downto 0);
  signal VGA_draw_count5 : std_logic_vector(4 downto 0);
  signal VGA_draw_count6 : std_logic_vector(4 downto 0);
  signal VGA_draw_count7 : std_logic_vector(4 downto 0);
  signal VGA_draw_count8 : std_logic_vector(4 downto 0);
  signal VGA_draw_count9 : std_logic_vector(4 downto 0);
  signal VGA_draw_count10 : std_logic_vector(4 downto 0);
  signal VGA_draw_count1 : std_logic_vector(4 downto 0);
  signal VGA_draw_count4 : std_logic_vector(4 downto 0);
  signal VGA_draw_count2 : std_logic_vector(4 downto 0);
  signal VGA_draw_count3 : std_logic_vector(4 downto 0);
  signal Collision_L1_range_state_out : std_logic_vector(1 downto 0);
  signal Collision_count_2_s : std_logic_vector(3 downto 0);
  signal Collision_count_1_s : std_logic_vector(3 downto 0);
  signal Collision_start_value_s : std_logic_vector(3 downto 0);
  signal Collision_L1_state : std_logic_vector(2 downto 0);
  signal Collision_L1_n_1, Collision_L1_n_2, Collision_L1_n_3, Collision_L1_n_4, Collision_L1_n_5 : std_logic;
  signal Collision_L1_n_6, Collision_L1_n_7, Collision_L1_n_8, Collision_L1_n_9, Collision_L1_n_10 : std_logic;
  signal Collision_L1_n_11, Collision_L1_n_12, Collision_L1_n_13, Collision_L1_n_14, Collision_L1_n_15 : std_logic;
  signal Collision_L1_n_16, Collision_L1_n_17, Collision_L1_n_18, Collision_L1_n_19, Collision_L1_n_20 : std_logic;
  signal Collision_L1_n_21, Collision_L1_n_22, Collision_L1_n_23, Collision_L1_n_24, Collision_L1_n_25 : std_logic;
  signal Collision_L1_n_26, Collision_L1_n_27, Collision_L1_n_28, Collision_L1_n_29, Collision_L1_n_30 : std_logic;
  signal Collision_L1_n_31, Collision_L1_n_32, Collision_L1_n_33, Collision_L1_n_34, Collision_L1_n_35 : std_logic;
  signal Collision_L1_n_36, Collision_L1_n_37, Collision_L1_n_38, Collision_L1_n_39, Collision_L1_n_40 : std_logic;
  signal Collision_L1_n_41, Collision_L1_n_42, Collision_L1_n_43, Collision_L1_n_44, Collision_L1_n_45 : std_logic;
  signal Collision_L1_n_46, Collision_L1_n_47, Collision_L1_n_48, Collision_L1_n_49, Collision_L1_n_50 : std_logic;
  signal Collision_L1_n_51, Collision_L1_n_52, Collision_L1_n_53, Collision_L1_n_54, Collision_L1_n_55 : std_logic;
  signal Collision_L1_n_56, Collision_L1_n_57, Collision_L1_n_58, Collision_L1_n_59, Collision_L1_n_60 : std_logic;
  signal Collision_L1_n_61, Collision_L1_n_62, Collision_L1_n_63, Collision_L1_n_64, Collision_L1_n_65 : std_logic;
  signal Collision_L1_n_66, Collision_L1_n_67, Collision_L1_n_68, Collision_L1_n_69, Collision_L1_n_70 : std_logic;
  signal Collision_L1_n_71, Collision_L1_n_72, Collision_L1_n_73, Collision_L1_n_74, Collision_L1_n_75 : std_logic;
  signal Collision_L1_n_76, Collision_L1_n_77, Collision_L1_n_78, Collision_L1_n_79, Collision_L1_n_80 : std_logic;
  signal Collision_L1_n_81, Collision_L1_n_82, Collision_L1_n_83, Collision_L1_n_84, Collision_L1_n_85 : std_logic;
  signal Collision_L1_n_86, Collision_L1_n_87, Collision_L1_n_88, Collision_L1_n_89, Collision_L1_n_90 : std_logic;
  signal Collision_L1_n_91, Collision_L1_n_92, Collision_L1_n_93, Collision_L1_n_94, Collision_L1_n_95 : std_logic;
  signal Collision_L1_n_96, Collision_L1_n_97, Collision_L1_n_98, Collision_L1_n_99, Collision_L1_n_100 : std_logic;
  signal Collision_L1_n_101, Collision_L1_n_102, Collision_L1_n_103, Collision_L1_n_104, Collision_L1_n_105 : std_logic;
  signal Collision_L1_n_106, Collision_L1_n_107, Collision_L1_n_108, Collision_L1_n_109, Collision_L1_n_110 : std_logic;
  signal Collision_L1_n_111, Collision_L1_n_112, Collision_L1_n_113, Collision_L1_n_114, Collision_L1_n_115 : std_logic;
  signal Collision_L1_n_116, Collision_L1_n_117, Collision_L1_n_118, Collision_L1_n_119, Collision_L1_n_120 : std_logic;
  signal Collision_L1_n_121, Collision_L1_n_122, Collision_L1_n_123, Collision_L1_n_124, Collision_L1_n_125 : std_logic;
  signal Collision_L1_n_126, Collision_L1_n_127, Collision_L1_n_128, Collision_L1_n_129, Collision_L1_n_130 : std_logic;
  signal Collision_L1_n_131, Collision_L1_n_132, Collision_L1_n_133, Collision_L1_n_134, Collision_L1_n_135 : std_logic;
  signal Collision_L1_n_136, Collision_L1_n_137, Collision_L1_n_138, Collision_L1_n_139, Collision_L1_n_140 : std_logic;
  signal Collision_L1_n_141, Collision_L1_n_142, Collision_L1_n_143, Collision_L1_n_144, Collision_L1_n_145 : std_logic;
  signal Collision_L1_n_146, Collision_L1_n_147, Collision_L1_n_148, Collision_L1_n_149, Collision_L1_n_150 : std_logic;
  signal Collision_L1_n_151, Collision_L1_n_152, Collision_L1_n_153, Collision_L1_n_154, Collision_L1_n_155 : std_logic;
  signal Collision_L1_n_156, Collision_L1_n_157, Collision_L1_n_158, Collision_L1_n_159, Collision_L1_n_160 : std_logic;
  signal Collision_L1_n_161, Collision_L1_n_162, Collision_L1_n_163, Collision_L1_n_164, Collision_L1_n_165 : std_logic;
  signal Collision_L1_n_166, Collision_L1_n_167, Collision_L1_n_168, Collision_L1_n_169, Collision_L1_n_170 : std_logic;
  signal Collision_L1_n_171, Collision_L1_n_172, Collision_L1_n_173, Collision_L1_n_174, Collision_L1_n_175 : std_logic;
  signal Collision_L1_n_176, Collision_L1_n_177, Collision_L1_n_178, Collision_L1_n_179, Collision_L1_n_180 : std_logic;
  signal Collision_L1_n_181, Collision_L1_n_182, Collision_L1_n_183, Collision_L1_n_184, Collision_L1_n_185 : std_logic;
  signal Collision_L1_n_186, Collision_L1_n_187, Collision_L1_n_188, Collision_L1_n_189, Collision_L1_n_190 : std_logic;
  signal Collision_L1_n_191, Collision_L1_n_192, Collision_L1_n_193, Collision_L1_n_194, Collision_L1_n_195 : std_logic;
  signal Collision_L1_n_196, Collision_L1_n_197, Collision_L1_n_198, Collision_L1_n_199, Collision_L1_n_200 : std_logic;
  signal Collision_L1_n_201, Collision_L1_n_202, Collision_L1_n_203, Collision_L1_n_204, Collision_L1_n_205 : std_logic;
  signal Collision_L1_n_206, Collision_L1_n_207, Collision_L1_n_208, Collision_L1_n_209, Collision_L1_n_210 : std_logic;
  signal Collision_L1_n_211, Collision_L1_n_212, Collision_L1_n_213, Collision_L1_n_214, Collision_L1_n_215 : std_logic;
  signal Collision_L1_n_216, Collision_L1_n_217, Collision_L1_n_218, Collision_L1_n_219, Collision_L1_n_220 : std_logic;
  signal Collision_L1_n_221, Collision_L1_n_222, Collision_L1_n_223, Collision_L1_n_224, Collision_L1_n_225 : std_logic;
  signal Collision_L1_n_226, Collision_L1_n_227, Collision_L1_n_228, Collision_L1_n_229, Collision_L1_n_230 : std_logic;
  signal Collision_L1_n_231, Collision_L1_n_232, Collision_L1_n_233, Collision_L1_n_234, Collision_L1_n_235 : std_logic;
  signal Collision_L1_n_236, Collision_L1_n_237, Collision_L1_n_238, Collision_L1_n_239, Collision_L1_n_240 : std_logic;
  signal Collision_L1_n_241, Collision_L1_n_242, Collision_L1_n_243, Collision_L1_n_244, Collision_L1_n_245 : std_logic;
  signal Collision_L1_n_246, Collision_L1_n_247, Collision_L1_n_248, Collision_L1_n_249, Collision_L1_n_250 : std_logic;
  signal Collision_L1_n_251, Collision_L1_n_252, Collision_L1_n_253, Collision_L1_n_254, Collision_L1_n_255 : std_logic;
  signal Collision_L1_n_256, Collision_L1_n_257, Collision_L1_n_258, Collision_L1_n_259, Collision_L1_n_260 : std_logic;
  signal Collision_L1_n_261, Collision_L1_n_262, Collision_L1_n_263, Collision_L1_n_264, Collision_L1_n_265 : std_logic;
  signal Collision_L1_n_266, Collision_L1_n_267, Collision_L1_n_268, Collision_L1_n_269, Collision_L1_n_270 : std_logic;
  signal Collision_L1_n_271, Collision_L1_n_272, Collision_L1_n_273, Collision_L1_n_274, Collision_L1_n_275 : std_logic;
  signal Collision_L1_n_276, Collision_L1_n_277, Collision_L1_n_278, Collision_L1_n_280, Collision_L1_n_281 : std_logic;
  signal Collision_L1_n_282, Collision_L1_n_283, Collision_L1_n_284, Collision_L1_n_285, Collision_L1_n_286 : std_logic;
  signal Collision_L1_n_287, Collision_L1_n_288, Collision_L1_n_289, Collision_L1_n_290, Collision_L1_n_291 : std_logic;
  signal Collision_L1_n_292, Collision_L1_n_293, Collision_L1_n_294, Collision_L1_n_295, Collision_L1_n_296 : std_logic;
  signal Collision_L1_n_297, Collision_L1_n_298, Collision_L1_n_299, Collision_L1_n_300, Collision_L1_n_301 : std_logic;
  signal Collision_L1_n_302, Collision_L1_n_303, Collision_L1_n_304, Collision_L1_n_305, Collision_L1_n_306 : std_logic;
  signal Collision_L1_n_307, Collision_L1_n_308, Collision_L1_n_309, Collision_L1_n_310, Collision_L1_n_311 : std_logic;
  signal Collision_L1_n_312, Collision_L1_n_313, Collision_L1_n_314, Collision_L1_n_315, Collision_L1_n_316 : std_logic;
  signal Collision_L1_n_317, Collision_L1_n_318, Collision_L1_n_319, Collision_L1_n_320, Collision_L1_n_321 : std_logic;
  signal Collision_L1_n_322, Collision_L1_n_323, Collision_L1_n_324, Collision_L1_n_325, Collision_L1_n_326 : std_logic;
  signal Collision_L1_n_327, Collision_L1_n_328, Collision_L1_n_329, Collision_L1_n_330, Collision_L1_n_331 : std_logic;
  signal Collision_L1_n_332, Collision_L1_n_333, Collision_L1_n_334, Collision_L1_n_335, Collision_L1_n_336 : std_logic;
  signal Collision_L1_n_337, Collision_L1_n_338, Collision_L1_n_339, Collision_L1_n_340, Collision_L1_n_341 : std_logic;
  signal Collision_L1_n_342, Collision_L1_n_343, Collision_L1_n_344, Collision_L1_n_345, Collision_L1_n_346 : std_logic;
  signal Collision_L1_n_347, Collision_L1_n_348, Collision_L1_n_349, Collision_L1_n_350, Collision_L1_n_351 : std_logic;
  signal Collision_L1_n_352, Collision_L1_n_353, Collision_L1_n_354, Collision_L1_n_355, Collision_L1_n_356 : std_logic;
  signal Collision_L1_n_357, Collision_L1_n_358, Collision_L1_n_359, Collision_L1_n_360, Collision_L1_n_361 : std_logic;
  signal Collision_L1_n_362, Collision_L1_n_363, Collision_L1_n_364, Collision_L1_n_365, Collision_L1_n_366 : std_logic;
  signal Collision_L1_n_367, Collision_L1_n_368, Collision_L1_n_369, Collision_L1_n_370, Collision_L1_n_371 : std_logic;
  signal Collision_L1_n_372, Collision_L1_n_373, Collision_L1_n_374, Collision_L1_n_375, Collision_L1_n_376 : std_logic;
  signal Collision_L1_n_377, Collision_L1_n_378, Collision_L1_n_380, Collision_L1_n_381, Collision_L1_n_382 : std_logic;
  signal Collision_L1_n_383, Collision_L1_n_385, Collision_L1_n_386, Collision_L1_n_387, Collision_L1_n_388 : std_logic;
  signal Collision_L1_n_389, Collision_L1_n_390, Collision_L1_n_391, Collision_L1_n_392, Collision_L1_n_393 : std_logic;
  signal Collision_L1_n_394, Collision_L1_n_395, Collision_L1_n_396, Collision_L1_n_399, Collision_L1_n_400 : std_logic;
  signal Collision_L1_n_401, Collision_L1_n_402, Collision_L1_n_403, Collision_L1_n_404, Collision_L1_n_405 : std_logic;
  signal Collision_L1_n_406, Collision_L1_n_407, Collision_L1_n_408, Collision_L1_n_409, Collision_L1_n_410 : std_logic;
  signal Collision_L1_n_411, Collision_L1_n_413, Collision_L1_n_415, Collision_L1_n_416, Collision_L1_n_417 : std_logic;
  signal Collision_L1_n_418, Collision_L1_n_419, Collision_L1_n_420, Collision_L1_n_421, Collision_L1_n_422 : std_logic;
  signal Collision_L1_n_423, Collision_L1_n_424, Collision_L1_n_425, Collision_L1_n_426, Collision_L1_n_427 : std_logic;
  signal Collision_L1_n_428, Collision_L1_n_429, Collision_L1_n_430, Collision_L1_n_431, Collision_L1_n_432 : std_logic;
  signal Collision_L1_n_433, Collision_L1_n_434, Collision_L1_n_435, Collision_L1_n_436, Collision_L1_n_437 : std_logic;
  signal Collision_L1_n_438, Collision_L1_n_439, Collision_L1_n_440, Collision_L1_n_441, Collision_L1_n_442 : std_logic;
  signal Collision_L1_n_443, Collision_L1_n_444, Collision_L1_n_445, Collision_L1_n_446, Collision_L1_n_447 : std_logic;
  signal Collision_L1_n_448, Collision_L1_n_449, Collision_L1_n_450, Collision_L1_n_451, Collision_L1_n_452 : std_logic;
  signal Collision_L1_n_453, Collision_L1_n_454, Collision_L1_n_455, Collision_L1_n_456, Collision_L1_n_457 : std_logic;
  signal Collision_L1_n_458, Collision_L1_n_459, Collision_L1_n_460, Collision_L1_n_461, Collision_L1_n_462 : std_logic;
  signal Collision_L1_n_463, Collision_L1_n_464, Collision_L1_n_465, Collision_L1_n_466, Collision_L1_n_467 : std_logic;
  signal Collision_L1_n_468, Collision_L1_n_469, Collision_L1_n_470, Collision_L1_n_471, Collision_L1_n_472 : std_logic;
  signal Collision_L1_n_473, Collision_L1_n_474, Collision_L1_n_475, Collision_L1_n_476, Collision_L1_n_479 : std_logic;
  signal Collision_L1_n_481, Collision_L1_n_482, Collision_L1_n_483, Collision_L1_n_484, Collision_L1_n_500 : std_logic;
  signal Collision_L1_n_501, Collision_L1_n_502, Collision_L1_n_503, Collision_L1_n_504, Collision_L1_n_505 : std_logic;
  signal Collision_L1_n_506, Collision_L1_n_509, Collision_L2_n_1, Collision_L2_n_2, Collision_L2_n_3 : std_logic;
  signal Collision_L2_n_4, Collision_L2_n_5, Collision_L2_n_6, Collision_L2_n_7, Collision_L2_n_8 : std_logic;
  signal Collision_L3_n_2, Collision_L3_n_3, Collision_L3_n_4, Collision_L3_n_5, Collision_L3_n_6 : std_logic;
  signal Collision_L3_n_7, Collision_L3_n_8, Collision_L3_n_9, Collision_L3_n_10, Collision_L3_n_11 : std_logic;
  signal Collision_L3_n_12, Collision_L3_n_13, Collision_enable_s, Collision_reset_2_s, Enemy_spawning_en11_n_0 : std_logic;
  signal Enemy_spawning_en11_n_1, Enemy_spawning_en11_n_2, Enemy_spawning_en11_n_3, Enemy_spawning_en21_n_0, Enemy_spawning_en21_n_1 : std_logic;
  signal Enemy_spawning_en21_n_2, Enemy_spawning_en21_n_3, Enemy_spawning_en31_n_0, Enemy_spawning_en31_n_1, Enemy_spawning_en31_n_2 : std_logic;
  signal Enemy_spawning_en31_n_3, Enemy_spawning_en41_n_0, Enemy_spawning_en41_n_1, Enemy_spawning_en41_n_2, Enemy_spawning_en41_n_3 : std_logic;
  signal Enemy_spawning_en51_n_0, Enemy_spawning_en51_n_1, Enemy_spawning_en51_n_2, Enemy_spawning_en51_n_3, Enemy_spawning_en61_n_0 : std_logic;
  signal Enemy_spawning_en61_n_1, Enemy_spawning_en61_n_2, Enemy_spawning_en61_n_3, Enemy_spawning_rngg_d1_n_0, Enemy_spawning_rngg_d2_n_0 : std_logic;
  signal Enemy_spawning_rngg_d3_n_0, Enemy_spawning_rngg_d4_n_0, Enemy_spawning_rngg_d5_n_0, Enemy_spawning_rngg_d6_n_0, Enemy_spawning_rngg_d7_n_0 : std_logic;
  signal Enemy_spawning_rngg_d8_n_0, Enemy_spawning_rngg_d9_n_0, Enemy_spawning_rngg_d10_n_0, Enemy_spawning_rngg_d11_n_0, Enemy_spawning_rngg_d12_n_0 : std_logic;
  signal Enemy_spawning_rngg_d13_n_0, Enemy_spawning_rngg_d14_n_0, Enemy_spawning_rngg_d15_n_0, Enemy_spawning_rngg_d16_n_0, Enemy_spawning_rngg_xor_input : std_logic;
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3 : std_logic;
  signal UNCONNECTED4, UNCONNECTED5, VGA_b1, VGA_b2, VGA_b3 : std_logic;
  signal VGA_b4, VGA_b5, VGA_b6, VGA_b7, VGA_b8 : std_logic;
  signal VGA_b9, VGA_b10, VGA_enable1, VGA_enable2, VGA_enable3 : std_logic;
  signal VGA_enable4, VGA_enable5, VGA_enable6, VGA_enable7, VGA_enable8 : std_logic;
  signal VGA_enable9, VGA_enable10, VGA_g1, VGA_g2, VGA_g3 : std_logic;
  signal VGA_g4, VGA_g5, VGA_g6, VGA_g7, VGA_g8 : std_logic;
  signal VGA_g9, VGA_g10, VGA_l01_n_2, VGA_l01_n_3, VGA_l01_n_4 : std_logic;
  signal VGA_l01_n_5, VGA_l01_n_6, VGA_l01_n_7, VGA_l01_n_8, VGA_l01_n_9 : std_logic;
  signal VGA_l01_n_10, VGA_l01_n_11, VGA_l01_n_12, VGA_l01_n_13, VGA_l01_n_14 : std_logic;
  signal VGA_l01_n_15, VGA_l01_n_16, VGA_l01_n_17, VGA_l01_n_18, VGA_l01_n_19 : std_logic;
  signal VGA_l01_n_20, VGA_l01_n_21, VGA_l01_n_22, VGA_l01_n_23, VGA_l01_n_24 : std_logic;
  signal VGA_l01_n_25, VGA_l01_n_26, VGA_l01_n_27, VGA_l01_n_28, VGA_l01_n_29 : std_logic;
  signal VGA_l01_n_30, VGA_l01_n_31, VGA_l01_n_32, VGA_l02_n_0, VGA_l02_n_1 : std_logic;
  signal VGA_l02_n_4, VGA_l02_n_5, VGA_l02_n_6, VGA_l02_n_7, VGA_l02_n_8 : std_logic;
  signal VGA_l02_n_9, VGA_l02_n_10, VGA_l02_n_11, VGA_l02_n_12, VGA_l02_n_13 : std_logic;
  signal VGA_l02_n_14, VGA_l02_n_15, VGA_l02_n_16, VGA_l02_n_17, VGA_l02_n_18 : std_logic;
  signal VGA_l02_n_19, VGA_l02_n_20, VGA_l02_n_21, VGA_l02_n_22, VGA_l02_n_23 : std_logic;
  signal VGA_l02_n_24, VGA_l02_n_25, VGA_l02_n_26, VGA_l02_n_27, VGA_l02_n_28 : std_logic;
  signal VGA_l02_n_29, VGA_l02_n_30, VGA_l02_n_31, VGA_l02_n_32, VGA_l02_n_33 : std_logic;
  signal VGA_l02_n_34, VGA_l02_n_35, VGA_l02_n_36, VGA_l02_n_37, VGA_l02_n_38 : std_logic;
  signal VGA_l02_n_39, VGA_l02_n_40, VGA_l03_n_2, VGA_l03_n_3, VGA_l03_n_4 : std_logic;
  signal VGA_l03_n_5, VGA_l03_n_6, VGA_l03_n_7, VGA_l03_n_8, VGA_l03_n_11 : std_logic;
  signal VGA_l03_n_12, VGA_l03_n_13, VGA_l03_n_35, VGA_l03_n_36, VGA_l06_n_0 : std_logic;
  signal VGA_l06_n_1, VGA_l06_n_2, VGA_l06_n_3, VGA_l06_n_4, VGA_l06_n_5 : std_logic;
  signal VGA_l06_n_6, VGA_l06_n_7, VGA_l06_n_8, VGA_l06_n_9, VGA_l06_n_10 : std_logic;
  signal VGA_l06_n_11, VGA_l06_n_12, VGA_l06_n_13, VGA_l06_n_14, VGA_l06_n_15 : std_logic;
  signal VGA_l06_n_16, VGA_l06_n_17, VGA_l06_n_18, VGA_l06_n_19, VGA_l06_n_20 : std_logic;
  signal VGA_l06_n_21, VGA_l06_n_22, VGA_l06_n_23, VGA_l06_n_24, VGA_l06_n_25 : std_logic;
  signal VGA_l06_n_26, VGA_l06_n_27, VGA_l06_n_28, VGA_l06_n_29, VGA_l06_n_30 : std_logic;
  signal VGA_l06_n_31, VGA_l06_n_32, VGA_l06_n_33, VGA_l06_n_34, VGA_l06_n_35 : std_logic;
  signal VGA_l06_n_36, VGA_l06_n_37, VGA_l06_n_38, VGA_l06_n_39, VGA_l06_n_40 : std_logic;
  signal VGA_l06_n_41, VGA_l06_n_42, VGA_l06_n_43, VGA_l06_n_44, VGA_l06_n_45 : std_logic;
  signal VGA_l06_n_46, VGA_l06_n_47, VGA_l06_n_48, VGA_l06_n_49, VGA_l06_n_50 : std_logic;
  signal VGA_l06_n_51, VGA_l06_n_52, VGA_l06_n_53, VGA_l06_n_54, VGA_l06_n_55 : std_logic;
  signal VGA_l06_n_56, VGA_l06_n_57, VGA_l06_n_58, VGA_l06_n_59, VGA_l06_n_60 : std_logic;
  signal VGA_l06_n_61, VGA_l06_n_62, VGA_l06_n_63, VGA_l06_n_64, VGA_l06_n_65 : std_logic;
  signal VGA_l06_n_66, VGA_l06_n_67, VGA_l06_n_68, VGA_l06_n_69, VGA_l06_n_70 : std_logic;
  signal VGA_l06_n_71, VGA_l06_n_72, VGA_l06_n_73, VGA_l06_n_74, VGA_l06_n_75 : std_logic;
  signal VGA_l06_n_76, VGA_l06_n_77, VGA_l06_n_78, VGA_l06_n_79, VGA_l06_n_80 : std_logic;
  signal VGA_l06_n_81, VGA_l06_n_82, VGA_l06_n_83, VGA_l06_n_84, VGA_l06_n_85 : std_logic;
  signal VGA_l06_n_86, VGA_l06_n_87, VGA_l06_n_88, VGA_l06_n_89, VGA_l06_n_90 : std_logic;
  signal VGA_l06_n_91, VGA_l06_n_92, VGA_l06_n_93, VGA_l06_n_94, VGA_l06_n_95 : std_logic;
  signal VGA_l06_n_96, VGA_l06_n_97, VGA_l06_n_98, VGA_l06_n_99, VGA_l06_n_100 : std_logic;
  signal VGA_l06_n_101, VGA_l06_n_102, VGA_l06_n_103, VGA_l06_n_104, VGA_l06_n_105 : std_logic;
  signal VGA_l06_n_106, VGA_l06_n_107, VGA_l06_n_108, VGA_l06_n_109, VGA_l06_n_110 : std_logic;
  signal VGA_l06_n_111, VGA_l06_n_112, VGA_l06_n_113, VGA_l06_n_114, VGA_l06_n_115 : std_logic;
  signal VGA_l06_n_116, VGA_l06_n_117, VGA_l06_n_118, VGA_l06_n_119, VGA_l06_n_120 : std_logic;
  signal VGA_l06_n_121, VGA_l06_n_122, VGA_l06_n_123, VGA_l06_n_124, VGA_l06_n_125 : std_logic;
  signal VGA_l06_n_126, VGA_l06_n_127, VGA_l06_n_128, VGA_l06_n_129, VGA_l06_n_130 : std_logic;
  signal VGA_l06_n_131, VGA_l06_n_132, VGA_l06_n_133, VGA_l06_n_134, VGA_l06_n_135 : std_logic;
  signal VGA_l06_n_136, VGA_l06_n_137, VGA_l06_n_138, VGA_l06_n_139, VGA_l06_n_140 : std_logic;
  signal VGA_l06_n_141, VGA_l06_n_142, VGA_l06_n_143, VGA_l06_n_144, VGA_l06_n_145 : std_logic;
  signal VGA_l06_n_146, VGA_l06_n_147, VGA_l06_n_148, VGA_l06_n_149, VGA_l06_n_150 : std_logic;
  signal VGA_l06_n_151, VGA_l06_n_152, VGA_l06_n_153, VGA_l06_n_154, VGA_l06_n_155 : std_logic;
  signal VGA_l06_n_156, VGA_l06_n_157, VGA_l06_n_158, VGA_l06_n_159, VGA_l06_n_160 : std_logic;
  signal VGA_l06_n_161, VGA_l06_n_162, VGA_l06_n_163, VGA_l06_n_164, VGA_l06_n_165 : std_logic;
  signal VGA_l06_n_166, VGA_l06_n_167, VGA_l06_n_168, VGA_l06_n_169, VGA_l06_n_170 : std_logic;
  signal VGA_l06_n_171, VGA_l06_n_172, VGA_l06_n_173, VGA_l06_n_174, VGA_l06_n_175 : std_logic;
  signal VGA_l06_n_176, VGA_l06_n_177, VGA_l06_n_178, VGA_l06_n_179, VGA_l06_n_180 : std_logic;
  signal VGA_l06_n_181, VGA_l06_n_182, VGA_l06_n_183, VGA_l06_n_184, VGA_l06_n_185 : std_logic;
  signal VGA_l06_n_186, VGA_l06_n_187, VGA_l06_n_188, VGA_l06_n_189, VGA_l06_n_190 : std_logic;
  signal VGA_l06_n_191, VGA_l06_n_192, VGA_l06_n_193, VGA_l06_n_194, VGA_l06_n_195 : std_logic;
  signal VGA_l06_n_196, VGA_l06_n_197, VGA_l06_n_198, VGA_l06_n_199, VGA_l06_n_200 : std_logic;
  signal VGA_l06_n_201, VGA_l06_n_202, VGA_l06_n_203, VGA_l06_n_204, VGA_l06_n_205 : std_logic;
  signal VGA_l06_n_206, VGA_l06_n_207, VGA_l06_n_208, VGA_l06_n_209, VGA_l06_n_210 : std_logic;
  signal VGA_l06_n_211, VGA_l06_n_212, VGA_l06_n_213, VGA_l06_n_214, VGA_l06_n_215 : std_logic;
  signal VGA_l06_n_216, VGA_l06_n_217, VGA_l06_n_218, VGA_l06_n_219, VGA_l06_n_220 : std_logic;
  signal VGA_l06_n_221, VGA_l06_n_222, VGA_l06_n_223, VGA_l06_n_224, VGA_l06_n_225 : std_logic;
  signal VGA_l06_n_226, VGA_l06_n_227, VGA_l06_n_228, VGA_l06_n_229, VGA_l06_n_230 : std_logic;
  signal VGA_l06_n_231, VGA_l06_n_232, VGA_l06_n_233, VGA_l06_n_234, VGA_l06_n_235 : std_logic;
  signal VGA_l06_n_236, VGA_l06_n_237, VGA_l06_n_238, VGA_l06_n_239, VGA_l06_n_240 : std_logic;
  signal VGA_l06_n_241, VGA_l06_n_242, VGA_l06_n_243, VGA_l06_n_244, VGA_l06_n_245 : std_logic;
  signal VGA_l06_n_246, VGA_l06_n_247, VGA_l06_n_248, VGA_l06_n_249, VGA_l06_n_250 : std_logic;
  signal VGA_l06_n_251, VGA_l06_n_252, VGA_l06_n_253, VGA_l06_n_254, VGA_l06_n_255 : std_logic;
  signal VGA_l06_n_256, VGA_l06_n_257, VGA_l06_n_258, VGA_l06_n_259, VGA_l06_n_260 : std_logic;
  signal VGA_l06_n_261, VGA_l06_n_262, VGA_l06_n_263, VGA_l06_n_264, VGA_l06_n_265 : std_logic;
  signal VGA_l06_n_266, VGA_l06_n_267, VGA_l06_n_268, VGA_l06_n_269, VGA_l06_n_270 : std_logic;
  signal VGA_l06_n_271, VGA_l06_n_272, VGA_l06_n_273, VGA_l06_n_274, VGA_l06_n_275 : std_logic;
  signal VGA_l06_n_276, VGA_l06_n_277, VGA_l06_n_278, VGA_l06_n_279, VGA_l06_n_280 : std_logic;
  signal VGA_l06_n_281, VGA_l06_n_282, VGA_l06_n_283, VGA_l06_n_284, VGA_l06_n_285 : std_logic;
  signal VGA_l06_n_286, VGA_l06_n_287, VGA_l06_n_288, VGA_l06_n_289, VGA_l06_n_290 : std_logic;
  signal VGA_l06_n_291, VGA_l06_n_292, VGA_l06_n_293, VGA_l06_n_294, VGA_l06_n_295 : std_logic;
  signal VGA_l06_n_296, VGA_l06_n_297, VGA_l06_n_298, VGA_l06_n_299, VGA_l06_n_300 : std_logic;
  signal VGA_l06_n_301, VGA_l06_n_302, VGA_l06_n_303, VGA_l06_n_304, VGA_l06_n_305 : std_logic;
  signal VGA_l06_n_306, VGA_l06_n_307, VGA_l06_n_308, VGA_l06_n_309, VGA_l06_n_310 : std_logic;
  signal VGA_l06_n_311, VGA_l06_n_312, VGA_l06_n_313, VGA_l06_n_314, VGA_l06_n_315 : std_logic;
  signal VGA_l06_n_316, VGA_l06_n_318, VGA_l06_n_319, VGA_l06_n_320, VGA_l06_n_322 : std_logic;
  signal VGA_l06_n_323, VGA_l041_n_0, VGA_l041_n_1, VGA_l041_n_2, VGA_l041_n_3 : std_logic;
  signal VGA_l041_n_4, VGA_l041_n_5, VGA_l041_n_6, VGA_l042_n_0, VGA_l042_n_1 : std_logic;
  signal VGA_l042_n_2, VGA_l042_n_3, VGA_l042_n_4, VGA_l042_n_5, VGA_l042_n_6 : std_logic;
  signal VGA_l043_n_0, VGA_l043_n_1, VGA_l043_n_2, VGA_l043_n_3, VGA_l043_n_4 : std_logic;
  signal VGA_l043_n_5, VGA_l043_n_6, VGA_l044_n_0, VGA_l044_n_1, VGA_l044_n_2 : std_logic;
  signal VGA_l044_n_3, VGA_l044_n_4, VGA_l044_n_5, VGA_l044_n_6, VGA_l044_n_7 : std_logic;
  signal VGA_l044_n_8, VGA_l044_n_9, VGA_l044_n_10, VGA_l044_n_11, VGA_l044_n_12 : std_logic;
  signal VGA_l045_n_0, VGA_l045_n_1, VGA_l045_n_2, VGA_l045_n_3, VGA_l045_n_4 : std_logic;
  signal VGA_l045_n_5, VGA_l045_n_6, VGA_l045_n_7, VGA_l045_n_8, VGA_l045_n_9 : std_logic;
  signal VGA_l045_n_10, VGA_l045_n_11, VGA_l045_n_12, VGA_l046_n_0, VGA_l046_n_1 : std_logic;
  signal VGA_l046_n_2, VGA_l046_n_3, VGA_l046_n_4, VGA_l046_n_5, VGA_l046_n_6 : std_logic;
  signal VGA_l046_n_7, VGA_l046_n_8, VGA_l046_n_9, VGA_l046_n_10, VGA_l046_n_11 : std_logic;
  signal VGA_l046_n_12, VGA_l047_n_0, VGA_l047_n_1, VGA_l047_n_2, VGA_l047_n_3 : std_logic;
  signal VGA_l047_n_4, VGA_l047_n_5, VGA_l047_n_6, VGA_l047_n_7, VGA_l047_n_8 : std_logic;
  signal VGA_l047_n_9, VGA_l047_n_10, VGA_l047_n_11, VGA_l047_n_12, VGA_l048_n_0 : std_logic;
  signal VGA_l048_n_1, VGA_l048_n_2, VGA_l048_n_3, VGA_l048_n_4, VGA_l048_n_5 : std_logic;
  signal VGA_l048_n_6, VGA_l048_n_7, VGA_l048_n_8, VGA_l048_n_9, VGA_l048_n_10 : std_logic;
  signal VGA_l048_n_11, VGA_l048_n_12, VGA_l049_n_0, VGA_l049_n_1, VGA_l049_n_2 : std_logic;
  signal VGA_l049_n_3, VGA_l049_n_4, VGA_l049_n_5, VGA_l049_n_6, VGA_l049_n_7 : std_logic;
  signal VGA_l049_n_8, VGA_l049_n_9, VGA_l049_n_10, VGA_l049_n_11, VGA_l049_n_12 : std_logic;
  signal VGA_l051_n_0, VGA_l051_n_1, VGA_l051_n_2, VGA_l051_n_3, VGA_l051_n_4 : std_logic;
  signal VGA_l051_n_5, VGA_l051_n_6, VGA_l051_n_7, VGA_l051_n_8, VGA_l051_n_9 : std_logic;
  signal VGA_l051_n_10, VGA_l051_n_11, VGA_l051_n_12, VGA_l051_n_13, VGA_l051_n_14 : std_logic;
  signal VGA_l051_n_15, VGA_l051_n_16, VGA_l051_n_17, VGA_l051_n_18, VGA_l051_n_19 : std_logic;
  signal VGA_l051_n_20, VGA_l051_n_21, VGA_l051_n_22, VGA_l051_n_23, VGA_l051_n_24 : std_logic;
  signal VGA_l051_n_25, VGA_l051_n_26, VGA_l051_n_27, VGA_l051_n_28, VGA_l051_n_29 : std_logic;
  signal VGA_l051_n_30, VGA_l051_n_31, VGA_l051_n_32, VGA_l051_n_33, VGA_l051_n_34 : std_logic;
  signal VGA_l051_n_35, VGA_l051_n_36, VGA_l051_n_37, VGA_l051_n_38, VGA_l051_n_39 : std_logic;
  signal VGA_l051_n_40, VGA_l051_n_41, VGA_l051_n_42, VGA_l051_n_43, VGA_l051_n_44 : std_logic;
  signal VGA_l051_n_45, VGA_l051_n_46, VGA_l051_n_47, VGA_l051_n_48, VGA_l051_n_49 : std_logic;
  signal VGA_l051_n_50, VGA_l051_n_51, VGA_l051_n_52, VGA_l051_n_53, VGA_l051_n_54 : std_logic;
  signal VGA_l051_n_55, VGA_l051_n_56, VGA_l051_n_57, VGA_l051_n_58, VGA_l051_n_59 : std_logic;
  signal VGA_l051_n_60, VGA_l051_n_61, VGA_l051_n_62, VGA_l051_n_63, VGA_l051_n_64 : std_logic;
  signal VGA_l051_n_65, VGA_l051_n_66, VGA_l051_n_67, VGA_l051_n_68, VGA_l051_n_69 : std_logic;
  signal VGA_l051_n_70, VGA_l051_n_71, VGA_l051_n_72, VGA_l051_n_73, VGA_l051_n_74 : std_logic;
  signal VGA_l051_n_75, VGA_l051_n_76, VGA_l051_n_77, VGA_l051_n_78, VGA_l051_n_79 : std_logic;
  signal VGA_l052_n_0, VGA_l052_n_1, VGA_l052_n_2, VGA_l052_n_3, VGA_l052_n_4 : std_logic;
  signal VGA_l052_n_5, VGA_l052_n_6, VGA_l052_n_7, VGA_l052_n_8, VGA_l052_n_9 : std_logic;
  signal VGA_l052_n_10, VGA_l052_n_11, VGA_l052_n_12, VGA_l052_n_13, VGA_l052_n_14 : std_logic;
  signal VGA_l052_n_15, VGA_l052_n_16, VGA_l052_n_17, VGA_l052_n_18, VGA_l052_n_19 : std_logic;
  signal VGA_l052_n_20, VGA_l052_n_21, VGA_l052_n_22, VGA_l052_n_23, VGA_l052_n_24 : std_logic;
  signal VGA_l052_n_25, VGA_l052_n_26, VGA_l052_n_27, VGA_l052_n_28, VGA_l052_n_29 : std_logic;
  signal VGA_l052_n_30, VGA_l052_n_31, VGA_l052_n_32, VGA_l052_n_33, VGA_l052_n_34 : std_logic;
  signal VGA_l052_n_35, VGA_l052_n_36, VGA_l052_n_37, VGA_l052_n_38, VGA_l052_n_39 : std_logic;
  signal VGA_l052_n_40, VGA_l052_n_41, VGA_l052_n_42, VGA_l052_n_43, VGA_l052_n_44 : std_logic;
  signal VGA_l052_n_45, VGA_l052_n_46, VGA_l052_n_47, VGA_l052_n_48, VGA_l052_n_49 : std_logic;
  signal VGA_l052_n_50, VGA_l052_n_51, VGA_l052_n_52, VGA_l052_n_53, VGA_l052_n_54 : std_logic;
  signal VGA_l052_n_55, VGA_l052_n_56, VGA_l052_n_57, VGA_l052_n_58, VGA_l052_n_59 : std_logic;
  signal VGA_l052_n_60, VGA_l052_n_61, VGA_l052_n_62, VGA_l052_n_63, VGA_l052_n_64 : std_logic;
  signal VGA_l052_n_65, VGA_l052_n_66, VGA_l052_n_67, VGA_l052_n_68, VGA_l052_n_69 : std_logic;
  signal VGA_l052_n_70, VGA_l052_n_71, VGA_l052_n_72, VGA_l052_n_73, VGA_l052_n_74 : std_logic;
  signal VGA_l052_n_75, VGA_l052_n_76, VGA_l052_n_77, VGA_l052_n_78, VGA_l052_n_79 : std_logic;
  signal VGA_l053_n_0, VGA_l053_n_1, VGA_l053_n_2, VGA_l053_n_3, VGA_l053_n_4 : std_logic;
  signal VGA_l053_n_5, VGA_l053_n_6, VGA_l053_n_7, VGA_l053_n_8, VGA_l053_n_9 : std_logic;
  signal VGA_l053_n_10, VGA_l053_n_11, VGA_l053_n_12, VGA_l053_n_13, VGA_l053_n_14 : std_logic;
  signal VGA_l053_n_15, VGA_l053_n_16, VGA_l053_n_17, VGA_l053_n_18, VGA_l053_n_19 : std_logic;
  signal VGA_l053_n_20, VGA_l053_n_21, VGA_l053_n_22, VGA_l053_n_23, VGA_l053_n_24 : std_logic;
  signal VGA_l053_n_25, VGA_l053_n_26, VGA_l053_n_27, VGA_l053_n_28, VGA_l053_n_29 : std_logic;
  signal VGA_l053_n_30, VGA_l053_n_31, VGA_l053_n_32, VGA_l053_n_33, VGA_l053_n_34 : std_logic;
  signal VGA_l053_n_35, VGA_l053_n_36, VGA_l053_n_37, VGA_l053_n_38, VGA_l053_n_39 : std_logic;
  signal VGA_l053_n_40, VGA_l053_n_41, VGA_l053_n_42, VGA_l053_n_43, VGA_l053_n_44 : std_logic;
  signal VGA_l053_n_45, VGA_l053_n_46, VGA_l053_n_47, VGA_l053_n_48, VGA_l053_n_49 : std_logic;
  signal VGA_l053_n_50, VGA_l053_n_51, VGA_l053_n_52, VGA_l053_n_53, VGA_l053_n_54 : std_logic;
  signal VGA_l053_n_55, VGA_l053_n_56, VGA_l053_n_57, VGA_l053_n_58, VGA_l053_n_59 : std_logic;
  signal VGA_l053_n_60, VGA_l053_n_61, VGA_l053_n_62, VGA_l053_n_63, VGA_l053_n_64 : std_logic;
  signal VGA_l053_n_65, VGA_l053_n_66, VGA_l053_n_67, VGA_l053_n_68, VGA_l053_n_69 : std_logic;
  signal VGA_l053_n_70, VGA_l053_n_71, VGA_l053_n_72, VGA_l053_n_73, VGA_l053_n_74 : std_logic;
  signal VGA_l053_n_75, VGA_l053_n_76, VGA_l053_n_77, VGA_l053_n_78, VGA_l053_n_79 : std_logic;
  signal VGA_l071_n_0, VGA_l071_n_1, VGA_l071_n_2, VGA_l071_n_3, VGA_l071_n_4 : std_logic;
  signal VGA_l071_n_5, VGA_l071_n_6, VGA_l071_n_7, VGA_l071_n_8, VGA_l071_n_9 : std_logic;
  signal VGA_l071_n_10, VGA_l071_n_11, VGA_l071_n_12, VGA_l071_n_13, VGA_l071_n_14 : std_logic;
  signal VGA_l071_n_15, VGA_l071_n_16, VGA_l071_n_17, VGA_l071_n_18, VGA_l071_n_19 : std_logic;
  signal VGA_l071_n_20, VGA_l071_n_21, VGA_l071_n_22, VGA_l071_n_23, VGA_l071_n_24 : std_logic;
  signal VGA_l071_n_25, VGA_l071_n_26, VGA_l071_n_27, VGA_l071_n_28, VGA_l071_n_29 : std_logic;
  signal VGA_l071_n_30, VGA_l071_n_31, VGA_l071_n_32, VGA_l071_n_33, VGA_l071_n_34 : std_logic;
  signal VGA_l071_n_35, VGA_l071_n_36, VGA_l071_n_37, VGA_l071_n_38, VGA_l071_n_39 : std_logic;
  signal VGA_l071_n_40, VGA_l071_n_41, VGA_l071_n_42, VGA_l071_n_43, VGA_l071_n_44 : std_logic;
  signal VGA_l071_n_45, VGA_l071_n_46, VGA_l071_n_47, VGA_l071_n_48, VGA_l071_n_49 : std_logic;
  signal VGA_l071_n_50, VGA_l071_n_51, VGA_l071_n_52, VGA_l071_n_53, VGA_l071_n_54 : std_logic;
  signal VGA_l071_n_55, VGA_l071_n_56, VGA_l071_n_57, VGA_l071_n_58, VGA_l071_n_59 : std_logic;
  signal VGA_l071_n_60, VGA_l071_n_61, VGA_l071_n_62, VGA_l071_n_63, VGA_l071_n_64 : std_logic;
  signal VGA_l071_n_65, VGA_l071_n_66, VGA_l071_n_67, VGA_l071_n_68, VGA_l071_n_69 : std_logic;
  signal VGA_l071_n_70, VGA_l071_n_71, VGA_l071_n_72, VGA_l071_n_73, VGA_l071_n_74 : std_logic;
  signal VGA_l071_n_75, VGA_l071_n_76, VGA_l071_n_77, VGA_l071_n_78, VGA_l071_n_79 : std_logic;
  signal VGA_l071_n_80, VGA_l071_n_81, VGA_l071_n_82, VGA_l071_n_83, VGA_l071_n_84 : std_logic;
  signal VGA_l071_n_85, VGA_l071_n_86, VGA_l071_n_87, VGA_l071_n_88, VGA_l071_n_89 : std_logic;
  signal VGA_l071_n_90, VGA_l071_n_91, VGA_l071_n_92, VGA_l071_n_93, VGA_l071_n_94 : std_logic;
  signal VGA_l071_n_95, VGA_l071_n_96, VGA_l071_n_97, VGA_l071_n_98, VGA_l071_n_99 : std_logic;
  signal VGA_l071_n_100, VGA_l071_n_101, VGA_l071_n_102, VGA_l071_n_103, VGA_l071_n_104 : std_logic;
  signal VGA_l071_n_105, VGA_l071_n_106, VGA_l071_n_107, VGA_l071_n_108, VGA_l071_n_109 : std_logic;
  signal VGA_l071_n_110, VGA_l071_n_111, VGA_l071_n_112, VGA_l071_n_113, VGA_l071_n_114 : std_logic;
  signal VGA_l071_n_115, VGA_l071_n_116, VGA_l071_n_117, VGA_l071_n_118, VGA_l071_n_119 : std_logic;
  signal VGA_l071_n_120, VGA_l071_n_121, VGA_l071_n_122, VGA_l071_n_123, VGA_l071_n_124 : std_logic;
  signal VGA_l071_n_125, VGA_l071_n_126, VGA_l071_n_127, VGA_l071_n_128, VGA_l071_n_129 : std_logic;
  signal VGA_l071_n_130, VGA_l071_n_131, VGA_l071_n_132, VGA_l071_n_133, VGA_l071_n_134 : std_logic;
  signal VGA_l071_n_135, VGA_l071_n_136, VGA_l071_n_137, VGA_l071_n_138, VGA_l071_n_139 : std_logic;
  signal VGA_l071_n_140, VGA_l071_n_141, VGA_l071_n_142, VGA_l071_n_143, VGA_l071_n_144 : std_logic;
  signal VGA_l071_n_145, VGA_l071_n_146, VGA_l071_n_147, VGA_l071_n_148, VGA_l071_n_149 : std_logic;
  signal VGA_l071_n_150, VGA_l071_n_151, VGA_l071_n_152, VGA_l071_n_153, VGA_l071_n_154 : std_logic;
  signal VGA_l071_n_155, VGA_l071_n_156, VGA_l071_n_157, VGA_l071_n_158, VGA_l071_n_159 : std_logic;
  signal VGA_l071_n_160, VGA_l071_n_161, VGA_l071_n_162, VGA_l071_n_163, VGA_l071_n_164 : std_logic;
  signal VGA_l071_n_165, VGA_l071_n_166, VGA_l071_n_167, VGA_l071_n_168, VGA_l071_n_169 : std_logic;
  signal VGA_l071_n_170, VGA_l071_n_171, VGA_l071_n_172, VGA_l071_n_173, VGA_l071_n_174 : std_logic;
  signal VGA_l071_n_175, VGA_l071_n_176, VGA_l071_n_177, VGA_l071_n_178, VGA_l071_n_179 : std_logic;
  signal VGA_l071_n_180, VGA_l071_n_181, VGA_l071_n_182, VGA_l071_n_183, VGA_l071_n_184 : std_logic;
  signal VGA_l071_n_185, VGA_l071_n_186, VGA_l071_n_187, VGA_l071_n_188, VGA_l071_n_189 : std_logic;
  signal VGA_l071_n_190, VGA_l071_n_191, VGA_l071_n_192, VGA_l071_n_193, VGA_l071_n_194 : std_logic;
  signal VGA_l071_n_195, VGA_l071_n_196, VGA_l071_n_197, VGA_l071_n_198, VGA_l071_n_199 : std_logic;
  signal VGA_l071_n_200, VGA_l071_n_201, VGA_l071_n_202, VGA_l071_n_203, VGA_l071_n_204 : std_logic;
  signal VGA_l071_n_205, VGA_l071_n_206, VGA_l071_n_207, VGA_l071_n_208, VGA_l071_n_209 : std_logic;
  signal VGA_l071_n_210, VGA_l071_n_211, VGA_l071_n_212, VGA_l071_n_213, VGA_l071_n_214 : std_logic;
  signal VGA_l071_n_215, VGA_l071_n_216, VGA_l071_n_217, VGA_l071_n_218, VGA_l071_n_219 : std_logic;
  signal VGA_l071_n_220, VGA_l071_n_221, VGA_l071_n_222, VGA_l071_n_223, VGA_l071_n_224 : std_logic;
  signal VGA_l071_n_225, VGA_l071_n_226, VGA_l071_n_227, VGA_l071_n_228, VGA_l071_n_229 : std_logic;
  signal VGA_l071_n_230, VGA_l071_n_231, VGA_l071_n_233, VGA_l071_n_235, VGA_l071_n_236 : std_logic;
  signal VGA_l071_n_237, VGA_l071_n_238, VGA_l071_n_239, VGA_l071_n_241, VGA_l071_n_242 : std_logic;
  signal VGA_l071_n_243, VGA_l072_n_0, VGA_l072_n_1, VGA_l072_n_2, VGA_l072_n_3 : std_logic;
  signal VGA_l072_n_4, VGA_l072_n_5, VGA_l072_n_6, VGA_l072_n_7, VGA_l072_n_8 : std_logic;
  signal VGA_l072_n_9, VGA_l072_n_10, VGA_l072_n_11, VGA_l072_n_12, VGA_l072_n_13 : std_logic;
  signal VGA_l072_n_14, VGA_l072_n_15, VGA_l072_n_16, VGA_l072_n_17, VGA_l072_n_18 : std_logic;
  signal VGA_l072_n_19, VGA_l072_n_20, VGA_l072_n_21, VGA_l072_n_22, VGA_l072_n_23 : std_logic;
  signal VGA_l072_n_24, VGA_l072_n_25, VGA_l072_n_26, VGA_l072_n_27, VGA_l072_n_28 : std_logic;
  signal VGA_l072_n_29, VGA_l072_n_30, VGA_l072_n_31, VGA_l072_n_32, VGA_l072_n_33 : std_logic;
  signal VGA_l072_n_34, VGA_l072_n_35, VGA_l072_n_36, VGA_l072_n_37, VGA_l072_n_38 : std_logic;
  signal VGA_l072_n_39, VGA_l072_n_40, VGA_l072_n_41, VGA_l072_n_42, VGA_l072_n_43 : std_logic;
  signal VGA_l072_n_44, VGA_l072_n_45, VGA_l072_n_46, VGA_l072_n_47, VGA_l072_n_48 : std_logic;
  signal VGA_l072_n_49, VGA_l072_n_50, VGA_l072_n_51, VGA_l072_n_52, VGA_l072_n_53 : std_logic;
  signal VGA_l072_n_54, VGA_l072_n_55, VGA_l072_n_56, VGA_l072_n_57, VGA_l072_n_58 : std_logic;
  signal VGA_l072_n_59, VGA_l072_n_60, VGA_l072_n_61, VGA_l072_n_62, VGA_l072_n_63 : std_logic;
  signal VGA_l072_n_64, VGA_l072_n_65, VGA_l072_n_66, VGA_l072_n_67, VGA_l072_n_68 : std_logic;
  signal VGA_l072_n_69, VGA_l072_n_70, VGA_l072_n_71, VGA_l072_n_72, VGA_l072_n_73 : std_logic;
  signal VGA_l072_n_74, VGA_l072_n_75, VGA_l072_n_76, VGA_l072_n_77, VGA_l072_n_78 : std_logic;
  signal VGA_l072_n_79, VGA_l072_n_80, VGA_l072_n_81, VGA_l072_n_82, VGA_l072_n_83 : std_logic;
  signal VGA_l072_n_84, VGA_l072_n_85, VGA_l072_n_86, VGA_l072_n_87, VGA_l072_n_88 : std_logic;
  signal VGA_l072_n_89, VGA_l072_n_90, VGA_l072_n_91, VGA_l072_n_92, VGA_l072_n_93 : std_logic;
  signal VGA_l072_n_94, VGA_l072_n_95, VGA_l072_n_96, VGA_l072_n_97, VGA_l072_n_98 : std_logic;
  signal VGA_l072_n_99, VGA_l072_n_100, VGA_l072_n_101, VGA_l072_n_102, VGA_l072_n_103 : std_logic;
  signal VGA_l072_n_104, VGA_l072_n_105, VGA_l072_n_106, VGA_l072_n_107, VGA_l072_n_108 : std_logic;
  signal VGA_l072_n_109, VGA_l072_n_110, VGA_l072_n_111, VGA_l072_n_112, VGA_l072_n_113 : std_logic;
  signal VGA_l072_n_114, VGA_l072_n_115, VGA_l072_n_116, VGA_l072_n_117, VGA_l072_n_118 : std_logic;
  signal VGA_l072_n_119, VGA_l072_n_120, VGA_l072_n_121, VGA_l072_n_122, VGA_l072_n_123 : std_logic;
  signal VGA_l072_n_124, VGA_l072_n_125, VGA_l072_n_126, VGA_l072_n_127, VGA_l072_n_128 : std_logic;
  signal VGA_l072_n_129, VGA_l072_n_130, VGA_l072_n_131, VGA_l072_n_132, VGA_l072_n_133 : std_logic;
  signal VGA_l072_n_134, VGA_l072_n_135, VGA_l072_n_136, VGA_l072_n_137, VGA_l072_n_138 : std_logic;
  signal VGA_l072_n_139, VGA_l072_n_140, VGA_l072_n_141, VGA_l072_n_142, VGA_l072_n_143 : std_logic;
  signal VGA_l072_n_144, VGA_l072_n_145, VGA_l072_n_146, VGA_l072_n_147, VGA_l072_n_148 : std_logic;
  signal VGA_l072_n_149, VGA_l072_n_150, VGA_l072_n_151, VGA_l072_n_152, VGA_l072_n_153 : std_logic;
  signal VGA_l072_n_154, VGA_l072_n_155, VGA_l072_n_156, VGA_l072_n_157, VGA_l072_n_158 : std_logic;
  signal VGA_l072_n_159, VGA_l072_n_160, VGA_l072_n_161, VGA_l072_n_162, VGA_l072_n_163 : std_logic;
  signal VGA_l072_n_164, VGA_l072_n_165, VGA_l072_n_166, VGA_l072_n_167, VGA_l072_n_168 : std_logic;
  signal VGA_l072_n_169, VGA_l072_n_170, VGA_l072_n_171, VGA_l072_n_172, VGA_l072_n_173 : std_logic;
  signal VGA_l072_n_174, VGA_l072_n_175, VGA_l072_n_176, VGA_l072_n_177, VGA_l072_n_178 : std_logic;
  signal VGA_l072_n_179, VGA_l072_n_180, VGA_l072_n_181, VGA_l072_n_182, VGA_l072_n_183 : std_logic;
  signal VGA_l072_n_184, VGA_l072_n_185, VGA_l072_n_186, VGA_l072_n_187, VGA_l072_n_188 : std_logic;
  signal VGA_l072_n_189, VGA_l072_n_190, VGA_l072_n_191, VGA_l072_n_192, VGA_l072_n_193 : std_logic;
  signal VGA_l072_n_194, VGA_l072_n_195, VGA_l072_n_196, VGA_l072_n_197, VGA_l072_n_198 : std_logic;
  signal VGA_l072_n_199, VGA_l072_n_200, VGA_l072_n_201, VGA_l072_n_202, VGA_l072_n_203 : std_logic;
  signal VGA_l072_n_204, VGA_l072_n_205, VGA_l072_n_206, VGA_l072_n_207, VGA_l072_n_208 : std_logic;
  signal VGA_l072_n_209, VGA_l072_n_210, VGA_l072_n_211, VGA_l072_n_212, VGA_l072_n_213 : std_logic;
  signal VGA_l072_n_214, VGA_l072_n_215, VGA_l072_n_216, VGA_l072_n_217, VGA_l072_n_218 : std_logic;
  signal VGA_l072_n_219, VGA_l072_n_220, VGA_l072_n_221, VGA_l072_n_222, VGA_l072_n_223 : std_logic;
  signal VGA_l072_n_224, VGA_l072_n_225, VGA_l072_n_226, VGA_l072_n_227, VGA_l072_n_228 : std_logic;
  signal VGA_l072_n_229, VGA_l072_n_230, VGA_l072_n_231, VGA_l072_n_233, VGA_l072_n_235 : std_logic;
  signal VGA_l072_n_236, VGA_l072_n_237, VGA_l072_n_238, VGA_l072_n_239, VGA_l072_n_241 : std_logic;
  signal VGA_l072_n_242, VGA_l072_n_243, VGA_l073_n_0, VGA_l073_n_1, VGA_l073_n_2 : std_logic;
  signal VGA_l073_n_3, VGA_l073_n_4, VGA_l073_n_5, VGA_l073_n_6, VGA_l073_n_7 : std_logic;
  signal VGA_l073_n_8, VGA_l073_n_9, VGA_l073_n_10, VGA_l073_n_11, VGA_l073_n_12 : std_logic;
  signal VGA_l073_n_13, VGA_l073_n_14, VGA_l073_n_15, VGA_l073_n_16, VGA_l073_n_17 : std_logic;
  signal VGA_l073_n_18, VGA_l073_n_19, VGA_l073_n_20, VGA_l073_n_21, VGA_l073_n_22 : std_logic;
  signal VGA_l073_n_23, VGA_l073_n_24, VGA_l073_n_25, VGA_l073_n_26, VGA_l073_n_27 : std_logic;
  signal VGA_l073_n_28, VGA_l073_n_29, VGA_l073_n_30, VGA_l073_n_31, VGA_l073_n_32 : std_logic;
  signal VGA_l073_n_33, VGA_l073_n_34, VGA_l073_n_35, VGA_l073_n_36, VGA_l073_n_37 : std_logic;
  signal VGA_l073_n_38, VGA_l073_n_39, VGA_l073_n_40, VGA_l073_n_41, VGA_l073_n_42 : std_logic;
  signal VGA_l073_n_43, VGA_l073_n_44, VGA_l073_n_45, VGA_l073_n_46, VGA_l073_n_47 : std_logic;
  signal VGA_l073_n_48, VGA_l073_n_49, VGA_l073_n_50, VGA_l073_n_51, VGA_l073_n_52 : std_logic;
  signal VGA_l073_n_53, VGA_l073_n_54, VGA_l073_n_55, VGA_l073_n_56, VGA_l073_n_57 : std_logic;
  signal VGA_l073_n_58, VGA_l073_n_59, VGA_l073_n_60, VGA_l073_n_61, VGA_l073_n_62 : std_logic;
  signal VGA_l073_n_63, VGA_l073_n_64, VGA_l073_n_65, VGA_l073_n_66, VGA_l073_n_67 : std_logic;
  signal VGA_l073_n_68, VGA_l073_n_69, VGA_l073_n_70, VGA_l073_n_71, VGA_l073_n_72 : std_logic;
  signal VGA_l073_n_73, VGA_l073_n_74, VGA_l073_n_75, VGA_l073_n_76, VGA_l073_n_77 : std_logic;
  signal VGA_l073_n_78, VGA_l073_n_79, VGA_l073_n_80, VGA_l073_n_81, VGA_l073_n_82 : std_logic;
  signal VGA_l073_n_83, VGA_l073_n_84, VGA_l073_n_85, VGA_l073_n_86, VGA_l073_n_87 : std_logic;
  signal VGA_l073_n_88, VGA_l073_n_89, VGA_l073_n_90, VGA_l073_n_91, VGA_l073_n_92 : std_logic;
  signal VGA_l073_n_93, VGA_l073_n_94, VGA_l073_n_95, VGA_l073_n_96, VGA_l073_n_97 : std_logic;
  signal VGA_l073_n_98, VGA_l073_n_99, VGA_l073_n_100, VGA_l073_n_101, VGA_l073_n_102 : std_logic;
  signal VGA_l073_n_103, VGA_l073_n_104, VGA_l073_n_105, VGA_l073_n_106, VGA_l073_n_107 : std_logic;
  signal VGA_l073_n_108, VGA_l073_n_109, VGA_l073_n_110, VGA_l073_n_111, VGA_l073_n_112 : std_logic;
  signal VGA_l073_n_113, VGA_l073_n_114, VGA_l073_n_115, VGA_l073_n_116, VGA_l073_n_117 : std_logic;
  signal VGA_l073_n_118, VGA_l073_n_119, VGA_l073_n_120, VGA_l073_n_121, VGA_l073_n_122 : std_logic;
  signal VGA_l073_n_123, VGA_l073_n_124, VGA_l073_n_125, VGA_l073_n_126, VGA_l073_n_127 : std_logic;
  signal VGA_l073_n_128, VGA_l073_n_129, VGA_l073_n_130, VGA_l073_n_131, VGA_l073_n_132 : std_logic;
  signal VGA_l073_n_133, VGA_l073_n_134, VGA_l073_n_135, VGA_l073_n_136, VGA_l073_n_137 : std_logic;
  signal VGA_l073_n_138, VGA_l073_n_139, VGA_l073_n_140, VGA_l073_n_141, VGA_l073_n_142 : std_logic;
  signal VGA_l073_n_143, VGA_l073_n_144, VGA_l073_n_145, VGA_l073_n_146, VGA_l073_n_147 : std_logic;
  signal VGA_l073_n_148, VGA_l073_n_149, VGA_l073_n_150, VGA_l073_n_151, VGA_l073_n_152 : std_logic;
  signal VGA_l073_n_153, VGA_l073_n_154, VGA_l073_n_155, VGA_l073_n_156, VGA_l073_n_157 : std_logic;
  signal VGA_l073_n_158, VGA_l073_n_159, VGA_l073_n_160, VGA_l073_n_161, VGA_l073_n_162 : std_logic;
  signal VGA_l073_n_163, VGA_l073_n_164, VGA_l073_n_165, VGA_l073_n_166, VGA_l073_n_167 : std_logic;
  signal VGA_l073_n_168, VGA_l073_n_169, VGA_l073_n_170, VGA_l073_n_171, VGA_l073_n_172 : std_logic;
  signal VGA_l073_n_173, VGA_l073_n_174, VGA_l073_n_175, VGA_l073_n_176, VGA_l073_n_177 : std_logic;
  signal VGA_l073_n_178, VGA_l073_n_179, VGA_l073_n_180, VGA_l073_n_181, VGA_l073_n_182 : std_logic;
  signal VGA_l073_n_183, VGA_l073_n_184, VGA_l073_n_185, VGA_l073_n_186, VGA_l073_n_187 : std_logic;
  signal VGA_l073_n_188, VGA_l073_n_189, VGA_l073_n_190, VGA_l073_n_191, VGA_l073_n_192 : std_logic;
  signal VGA_l073_n_193, VGA_l073_n_194, VGA_l073_n_195, VGA_l073_n_196, VGA_l073_n_197 : std_logic;
  signal VGA_l073_n_198, VGA_l073_n_199, VGA_l073_n_200, VGA_l073_n_201, VGA_l073_n_202 : std_logic;
  signal VGA_l073_n_203, VGA_l073_n_204, VGA_l073_n_205, VGA_l073_n_206, VGA_l073_n_207 : std_logic;
  signal VGA_l073_n_208, VGA_l073_n_209, VGA_l073_n_210, VGA_l073_n_211, VGA_l073_n_212 : std_logic;
  signal VGA_l073_n_213, VGA_l073_n_214, VGA_l073_n_215, VGA_l073_n_216, VGA_l073_n_217 : std_logic;
  signal VGA_l073_n_218, VGA_l073_n_219, VGA_l073_n_220, VGA_l073_n_221, VGA_l073_n_222 : std_logic;
  signal VGA_l073_n_223, VGA_l073_n_224, VGA_l073_n_225, VGA_l073_n_226, VGA_l073_n_227 : std_logic;
  signal VGA_l073_n_228, VGA_l073_n_229, VGA_l073_n_230, VGA_l073_n_231, VGA_l073_n_233 : std_logic;
  signal VGA_l073_n_235, VGA_l073_n_236, VGA_l073_n_237, VGA_l073_n_238, VGA_l073_n_239 : std_logic;
  signal VGA_l073_n_241, VGA_l073_n_242, VGA_l073_n_243, VGA_l074_n_0, VGA_l074_n_1 : std_logic;
  signal VGA_l074_n_2, VGA_l074_n_3, VGA_l074_n_4, VGA_l074_n_5, VGA_l074_n_6 : std_logic;
  signal VGA_l074_n_7, VGA_l074_n_8, VGA_l074_n_9, VGA_l074_n_10, VGA_l074_n_11 : std_logic;
  signal VGA_l074_n_12, VGA_l074_n_13, VGA_l074_n_14, VGA_l074_n_15, VGA_l074_n_16 : std_logic;
  signal VGA_l074_n_17, VGA_l074_n_18, VGA_l074_n_19, VGA_l074_n_20, VGA_l074_n_21 : std_logic;
  signal VGA_l074_n_22, VGA_l074_n_23, VGA_l074_n_24, VGA_l074_n_25, VGA_l074_n_26 : std_logic;
  signal VGA_l074_n_27, VGA_l074_n_28, VGA_l074_n_29, VGA_l074_n_30, VGA_l074_n_31 : std_logic;
  signal VGA_l074_n_32, VGA_l074_n_33, VGA_l074_n_34, VGA_l074_n_35, VGA_l074_n_36 : std_logic;
  signal VGA_l074_n_37, VGA_l074_n_38, VGA_l074_n_39, VGA_l074_n_40, VGA_l074_n_41 : std_logic;
  signal VGA_l074_n_42, VGA_l074_n_43, VGA_l074_n_44, VGA_l074_n_45, VGA_l074_n_46 : std_logic;
  signal VGA_l074_n_47, VGA_l074_n_48, VGA_l074_n_49, VGA_l074_n_50, VGA_l074_n_51 : std_logic;
  signal VGA_l074_n_52, VGA_l074_n_53, VGA_l074_n_54, VGA_l074_n_55, VGA_l074_n_56 : std_logic;
  signal VGA_l074_n_57, VGA_l074_n_58, VGA_l074_n_59, VGA_l074_n_60, VGA_l074_n_61 : std_logic;
  signal VGA_l074_n_62, VGA_l074_n_63, VGA_l074_n_64, VGA_l074_n_65, VGA_l074_n_66 : std_logic;
  signal VGA_l074_n_67, VGA_l074_n_68, VGA_l074_n_69, VGA_l074_n_70, VGA_l074_n_71 : std_logic;
  signal VGA_l074_n_72, VGA_l074_n_73, VGA_l074_n_74, VGA_l074_n_75, VGA_l074_n_76 : std_logic;
  signal VGA_l074_n_77, VGA_l074_n_78, VGA_l074_n_79, VGA_l074_n_80, VGA_l074_n_81 : std_logic;
  signal VGA_l074_n_82, VGA_l074_n_83, VGA_l074_n_84, VGA_l074_n_85, VGA_l074_n_86 : std_logic;
  signal VGA_l074_n_87, VGA_l074_n_88, VGA_l074_n_89, VGA_l074_n_90, VGA_l074_n_91 : std_logic;
  signal VGA_l074_n_92, VGA_l074_n_93, VGA_l074_n_94, VGA_l074_n_95, VGA_l074_n_96 : std_logic;
  signal VGA_l074_n_97, VGA_l074_n_98, VGA_l074_n_99, VGA_l074_n_100, VGA_l074_n_101 : std_logic;
  signal VGA_l074_n_102, VGA_l074_n_103, VGA_l074_n_104, VGA_l074_n_105, VGA_l074_n_106 : std_logic;
  signal VGA_l074_n_107, VGA_l074_n_108, VGA_l074_n_109, VGA_l074_n_110, VGA_l074_n_111 : std_logic;
  signal VGA_l074_n_112, VGA_l074_n_113, VGA_l074_n_114, VGA_l074_n_115, VGA_l074_n_116 : std_logic;
  signal VGA_l074_n_117, VGA_l074_n_118, VGA_l074_n_119, VGA_l074_n_120, VGA_l074_n_121 : std_logic;
  signal VGA_l074_n_122, VGA_l074_n_123, VGA_l074_n_124, VGA_l074_n_125, VGA_l074_n_126 : std_logic;
  signal VGA_l074_n_127, VGA_l074_n_128, VGA_l074_n_129, VGA_l074_n_130, VGA_l074_n_131 : std_logic;
  signal VGA_l074_n_132, VGA_l074_n_133, VGA_l074_n_134, VGA_l074_n_135, VGA_l074_n_136 : std_logic;
  signal VGA_l074_n_137, VGA_l074_n_138, VGA_l074_n_139, VGA_l074_n_140, VGA_l074_n_141 : std_logic;
  signal VGA_l074_n_142, VGA_l074_n_143, VGA_l074_n_144, VGA_l074_n_145, VGA_l074_n_146 : std_logic;
  signal VGA_l074_n_147, VGA_l074_n_148, VGA_l074_n_149, VGA_l074_n_150, VGA_l074_n_151 : std_logic;
  signal VGA_l074_n_152, VGA_l074_n_153, VGA_l074_n_154, VGA_l074_n_155, VGA_l074_n_156 : std_logic;
  signal VGA_l074_n_157, VGA_l074_n_158, VGA_l074_n_159, VGA_l074_n_160, VGA_l074_n_161 : std_logic;
  signal VGA_l074_n_162, VGA_l074_n_163, VGA_l074_n_164, VGA_l074_n_165, VGA_l074_n_166 : std_logic;
  signal VGA_l074_n_167, VGA_l074_n_168, VGA_l074_n_169, VGA_l074_n_170, VGA_l074_n_171 : std_logic;
  signal VGA_l074_n_172, VGA_l074_n_173, VGA_l074_n_174, VGA_l074_n_175, VGA_l074_n_176 : std_logic;
  signal VGA_l074_n_177, VGA_l074_n_178, VGA_l074_n_179, VGA_l074_n_180, VGA_l074_n_181 : std_logic;
  signal VGA_l074_n_182, VGA_l074_n_183, VGA_l074_n_184, VGA_l074_n_185, VGA_l074_n_186 : std_logic;
  signal VGA_l074_n_187, VGA_l074_n_188, VGA_l074_n_189, VGA_l074_n_190, VGA_l074_n_191 : std_logic;
  signal VGA_l074_n_192, VGA_l074_n_193, VGA_l074_n_194, VGA_l074_n_195, VGA_l074_n_196 : std_logic;
  signal VGA_l074_n_197, VGA_l074_n_198, VGA_l074_n_199, VGA_l074_n_200, VGA_l074_n_201 : std_logic;
  signal VGA_l074_n_202, VGA_l074_n_203, VGA_l074_n_204, VGA_l074_n_205, VGA_l074_n_206 : std_logic;
  signal VGA_l074_n_207, VGA_l074_n_208, VGA_l074_n_209, VGA_l074_n_210, VGA_l074_n_211 : std_logic;
  signal VGA_l074_n_212, VGA_l074_n_213, VGA_l074_n_214, VGA_l074_n_215, VGA_l074_n_216 : std_logic;
  signal VGA_l074_n_217, VGA_l074_n_218, VGA_l074_n_219, VGA_l074_n_220, VGA_l074_n_221 : std_logic;
  signal VGA_l074_n_222, VGA_l074_n_223, VGA_l074_n_224, VGA_l074_n_225, VGA_l074_n_226 : std_logic;
  signal VGA_l074_n_227, VGA_l074_n_228, VGA_l074_n_229, VGA_l074_n_230, VGA_l074_n_231 : std_logic;
  signal VGA_l074_n_233, VGA_l074_n_235, VGA_l074_n_236, VGA_l074_n_237, VGA_l074_n_238 : std_logic;
  signal VGA_l074_n_239, VGA_l074_n_241, VGA_l074_n_242, VGA_l074_n_243, VGA_l075_n_0 : std_logic;
  signal VGA_l075_n_1, VGA_l075_n_2, VGA_l075_n_3, VGA_l075_n_4, VGA_l075_n_5 : std_logic;
  signal VGA_l075_n_6, VGA_l075_n_7, VGA_l075_n_8, VGA_l075_n_9, VGA_l075_n_10 : std_logic;
  signal VGA_l075_n_11, VGA_l075_n_12, VGA_l075_n_13, VGA_l075_n_14, VGA_l075_n_15 : std_logic;
  signal VGA_l075_n_16, VGA_l075_n_17, VGA_l075_n_18, VGA_l075_n_19, VGA_l075_n_20 : std_logic;
  signal VGA_l075_n_21, VGA_l075_n_22, VGA_l075_n_23, VGA_l075_n_24, VGA_l075_n_25 : std_logic;
  signal VGA_l075_n_26, VGA_l075_n_27, VGA_l075_n_28, VGA_l075_n_29, VGA_l075_n_30 : std_logic;
  signal VGA_l075_n_31, VGA_l075_n_32, VGA_l075_n_33, VGA_l075_n_34, VGA_l075_n_35 : std_logic;
  signal VGA_l075_n_36, VGA_l075_n_37, VGA_l075_n_38, VGA_l075_n_39, VGA_l075_n_40 : std_logic;
  signal VGA_l075_n_41, VGA_l075_n_42, VGA_l075_n_43, VGA_l075_n_44, VGA_l075_n_45 : std_logic;
  signal VGA_l075_n_46, VGA_l075_n_47, VGA_l075_n_48, VGA_l075_n_49, VGA_l075_n_50 : std_logic;
  signal VGA_l075_n_51, VGA_l075_n_52, VGA_l075_n_53, VGA_l075_n_54, VGA_l075_n_55 : std_logic;
  signal VGA_l075_n_56, VGA_l075_n_57, VGA_l075_n_58, VGA_l075_n_59, VGA_l075_n_60 : std_logic;
  signal VGA_l075_n_61, VGA_l075_n_62, VGA_l075_n_63, VGA_l075_n_64, VGA_l075_n_65 : std_logic;
  signal VGA_l075_n_66, VGA_l075_n_67, VGA_l075_n_68, VGA_l075_n_69, VGA_l075_n_70 : std_logic;
  signal VGA_l075_n_71, VGA_l075_n_72, VGA_l075_n_73, VGA_l075_n_74, VGA_l075_n_75 : std_logic;
  signal VGA_l075_n_76, VGA_l075_n_77, VGA_l075_n_78, VGA_l075_n_79, VGA_l075_n_80 : std_logic;
  signal VGA_l075_n_81, VGA_l075_n_82, VGA_l075_n_83, VGA_l075_n_84, VGA_l075_n_85 : std_logic;
  signal VGA_l075_n_86, VGA_l075_n_87, VGA_l075_n_88, VGA_l075_n_89, VGA_l075_n_90 : std_logic;
  signal VGA_l075_n_91, VGA_l075_n_92, VGA_l075_n_93, VGA_l075_n_94, VGA_l075_n_95 : std_logic;
  signal VGA_l075_n_96, VGA_l075_n_97, VGA_l075_n_98, VGA_l075_n_99, VGA_l075_n_100 : std_logic;
  signal VGA_l075_n_101, VGA_l075_n_102, VGA_l075_n_103, VGA_l075_n_104, VGA_l075_n_105 : std_logic;
  signal VGA_l075_n_106, VGA_l075_n_107, VGA_l075_n_108, VGA_l075_n_109, VGA_l075_n_110 : std_logic;
  signal VGA_l075_n_111, VGA_l075_n_112, VGA_l075_n_113, VGA_l075_n_114, VGA_l075_n_115 : std_logic;
  signal VGA_l075_n_116, VGA_l075_n_117, VGA_l075_n_118, VGA_l075_n_119, VGA_l075_n_120 : std_logic;
  signal VGA_l075_n_121, VGA_l075_n_122, VGA_l075_n_123, VGA_l075_n_124, VGA_l075_n_125 : std_logic;
  signal VGA_l075_n_126, VGA_l075_n_127, VGA_l075_n_128, VGA_l075_n_129, VGA_l075_n_130 : std_logic;
  signal VGA_l075_n_131, VGA_l075_n_132, VGA_l075_n_133, VGA_l075_n_134, VGA_l075_n_135 : std_logic;
  signal VGA_l075_n_136, VGA_l075_n_137, VGA_l075_n_138, VGA_l075_n_139, VGA_l075_n_140 : std_logic;
  signal VGA_l075_n_141, VGA_l075_n_142, VGA_l075_n_143, VGA_l075_n_144, VGA_l075_n_145 : std_logic;
  signal VGA_l075_n_146, VGA_l075_n_147, VGA_l075_n_148, VGA_l075_n_149, VGA_l075_n_150 : std_logic;
  signal VGA_l075_n_151, VGA_l075_n_152, VGA_l075_n_153, VGA_l075_n_154, VGA_l075_n_155 : std_logic;
  signal VGA_l075_n_156, VGA_l075_n_157, VGA_l075_n_158, VGA_l075_n_159, VGA_l075_n_160 : std_logic;
  signal VGA_l075_n_161, VGA_l075_n_162, VGA_l075_n_163, VGA_l075_n_164, VGA_l075_n_165 : std_logic;
  signal VGA_l075_n_166, VGA_l075_n_167, VGA_l075_n_168, VGA_l075_n_169, VGA_l075_n_170 : std_logic;
  signal VGA_l075_n_171, VGA_l075_n_172, VGA_l075_n_173, VGA_l075_n_174, VGA_l075_n_175 : std_logic;
  signal VGA_l075_n_176, VGA_l075_n_177, VGA_l075_n_178, VGA_l075_n_179, VGA_l075_n_180 : std_logic;
  signal VGA_l075_n_181, VGA_l075_n_182, VGA_l075_n_183, VGA_l075_n_184, VGA_l075_n_185 : std_logic;
  signal VGA_l075_n_186, VGA_l075_n_187, VGA_l075_n_188, VGA_l075_n_189, VGA_l075_n_190 : std_logic;
  signal VGA_l075_n_191, VGA_l075_n_192, VGA_l075_n_193, VGA_l075_n_194, VGA_l075_n_195 : std_logic;
  signal VGA_l075_n_196, VGA_l075_n_197, VGA_l075_n_198, VGA_l075_n_199, VGA_l075_n_200 : std_logic;
  signal VGA_l075_n_201, VGA_l075_n_202, VGA_l075_n_203, VGA_l075_n_204, VGA_l075_n_205 : std_logic;
  signal VGA_l075_n_206, VGA_l075_n_207, VGA_l075_n_208, VGA_l075_n_209, VGA_l075_n_210 : std_logic;
  signal VGA_l075_n_211, VGA_l075_n_212, VGA_l075_n_213, VGA_l075_n_214, VGA_l075_n_215 : std_logic;
  signal VGA_l075_n_216, VGA_l075_n_217, VGA_l075_n_218, VGA_l075_n_219, VGA_l075_n_220 : std_logic;
  signal VGA_l075_n_221, VGA_l075_n_222, VGA_l075_n_223, VGA_l075_n_224, VGA_l075_n_225 : std_logic;
  signal VGA_l075_n_226, VGA_l075_n_227, VGA_l075_n_228, VGA_l075_n_229, VGA_l075_n_230 : std_logic;
  signal VGA_l075_n_231, VGA_l075_n_233, VGA_l075_n_235, VGA_l075_n_236, VGA_l075_n_237 : std_logic;
  signal VGA_l075_n_238, VGA_l075_n_239, VGA_l075_n_241, VGA_l075_n_242, VGA_l075_n_243 : std_logic;
  signal VGA_l076_n_0, VGA_l076_n_1, VGA_l076_n_2, VGA_l076_n_3, VGA_l076_n_4 : std_logic;
  signal VGA_l076_n_5, VGA_l076_n_6, VGA_l076_n_7, VGA_l076_n_8, VGA_l076_n_9 : std_logic;
  signal VGA_l076_n_10, VGA_l076_n_11, VGA_l076_n_12, VGA_l076_n_13, VGA_l076_n_14 : std_logic;
  signal VGA_l076_n_15, VGA_l076_n_16, VGA_l076_n_17, VGA_l076_n_18, VGA_l076_n_19 : std_logic;
  signal VGA_l076_n_20, VGA_l076_n_21, VGA_l076_n_22, VGA_l076_n_23, VGA_l076_n_24 : std_logic;
  signal VGA_l076_n_25, VGA_l076_n_26, VGA_l076_n_27, VGA_l076_n_28, VGA_l076_n_29 : std_logic;
  signal VGA_l076_n_30, VGA_l076_n_31, VGA_l076_n_32, VGA_l076_n_33, VGA_l076_n_34 : std_logic;
  signal VGA_l076_n_35, VGA_l076_n_36, VGA_l076_n_37, VGA_l076_n_38, VGA_l076_n_39 : std_logic;
  signal VGA_l076_n_40, VGA_l076_n_41, VGA_l076_n_42, VGA_l076_n_43, VGA_l076_n_44 : std_logic;
  signal VGA_l076_n_45, VGA_l076_n_46, VGA_l076_n_47, VGA_l076_n_48, VGA_l076_n_49 : std_logic;
  signal VGA_l076_n_50, VGA_l076_n_51, VGA_l076_n_52, VGA_l076_n_53, VGA_l076_n_54 : std_logic;
  signal VGA_l076_n_55, VGA_l076_n_56, VGA_l076_n_57, VGA_l076_n_58, VGA_l076_n_59 : std_logic;
  signal VGA_l076_n_60, VGA_l076_n_61, VGA_l076_n_62, VGA_l076_n_63, VGA_l076_n_64 : std_logic;
  signal VGA_l076_n_65, VGA_l076_n_66, VGA_l076_n_67, VGA_l076_n_68, VGA_l076_n_69 : std_logic;
  signal VGA_l076_n_70, VGA_l076_n_71, VGA_l076_n_72, VGA_l076_n_73, VGA_l076_n_74 : std_logic;
  signal VGA_l076_n_75, VGA_l076_n_76, VGA_l076_n_77, VGA_l076_n_78, VGA_l076_n_79 : std_logic;
  signal VGA_l076_n_80, VGA_l076_n_81, VGA_l076_n_82, VGA_l076_n_83, VGA_l076_n_84 : std_logic;
  signal VGA_l076_n_85, VGA_l076_n_86, VGA_l076_n_87, VGA_l076_n_88, VGA_l076_n_89 : std_logic;
  signal VGA_l076_n_90, VGA_l076_n_91, VGA_l076_n_92, VGA_l076_n_93, VGA_l076_n_94 : std_logic;
  signal VGA_l076_n_95, VGA_l076_n_96, VGA_l076_n_97, VGA_l076_n_98, VGA_l076_n_99 : std_logic;
  signal VGA_l076_n_100, VGA_l076_n_101, VGA_l076_n_102, VGA_l076_n_103, VGA_l076_n_104 : std_logic;
  signal VGA_l076_n_105, VGA_l076_n_106, VGA_l076_n_107, VGA_l076_n_108, VGA_l076_n_109 : std_logic;
  signal VGA_l076_n_110, VGA_l076_n_111, VGA_l076_n_112, VGA_l076_n_113, VGA_l076_n_114 : std_logic;
  signal VGA_l076_n_115, VGA_l076_n_116, VGA_l076_n_117, VGA_l076_n_118, VGA_l076_n_119 : std_logic;
  signal VGA_l076_n_120, VGA_l076_n_121, VGA_l076_n_122, VGA_l076_n_123, VGA_l076_n_124 : std_logic;
  signal VGA_l076_n_125, VGA_l076_n_126, VGA_l076_n_127, VGA_l076_n_128, VGA_l076_n_129 : std_logic;
  signal VGA_l076_n_130, VGA_l076_n_131, VGA_l076_n_132, VGA_l076_n_133, VGA_l076_n_134 : std_logic;
  signal VGA_l076_n_135, VGA_l076_n_136, VGA_l076_n_137, VGA_l076_n_138, VGA_l076_n_139 : std_logic;
  signal VGA_l076_n_140, VGA_l076_n_141, VGA_l076_n_142, VGA_l076_n_143, VGA_l076_n_144 : std_logic;
  signal VGA_l076_n_145, VGA_l076_n_146, VGA_l076_n_147, VGA_l076_n_148, VGA_l076_n_149 : std_logic;
  signal VGA_l076_n_150, VGA_l076_n_151, VGA_l076_n_152, VGA_l076_n_153, VGA_l076_n_154 : std_logic;
  signal VGA_l076_n_155, VGA_l076_n_156, VGA_l076_n_157, VGA_l076_n_158, VGA_l076_n_159 : std_logic;
  signal VGA_l076_n_160, VGA_l076_n_161, VGA_l076_n_162, VGA_l076_n_163, VGA_l076_n_164 : std_logic;
  signal VGA_l076_n_165, VGA_l076_n_166, VGA_l076_n_167, VGA_l076_n_168, VGA_l076_n_169 : std_logic;
  signal VGA_l076_n_170, VGA_l076_n_171, VGA_l076_n_172, VGA_l076_n_173, VGA_l076_n_174 : std_logic;
  signal VGA_l076_n_175, VGA_l076_n_176, VGA_l076_n_177, VGA_l076_n_178, VGA_l076_n_179 : std_logic;
  signal VGA_l076_n_180, VGA_l076_n_181, VGA_l076_n_182, VGA_l076_n_183, VGA_l076_n_184 : std_logic;
  signal VGA_l076_n_185, VGA_l076_n_186, VGA_l076_n_187, VGA_l076_n_188, VGA_l076_n_189 : std_logic;
  signal VGA_l076_n_190, VGA_l076_n_191, VGA_l076_n_192, VGA_l076_n_193, VGA_l076_n_194 : std_logic;
  signal VGA_l076_n_195, VGA_l076_n_196, VGA_l076_n_197, VGA_l076_n_198, VGA_l076_n_199 : std_logic;
  signal VGA_l076_n_200, VGA_l076_n_201, VGA_l076_n_202, VGA_l076_n_203, VGA_l076_n_204 : std_logic;
  signal VGA_l076_n_205, VGA_l076_n_206, VGA_l076_n_207, VGA_l076_n_208, VGA_l076_n_209 : std_logic;
  signal VGA_l076_n_210, VGA_l076_n_211, VGA_l076_n_212, VGA_l076_n_213, VGA_l076_n_214 : std_logic;
  signal VGA_l076_n_215, VGA_l076_n_216, VGA_l076_n_217, VGA_l076_n_218, VGA_l076_n_219 : std_logic;
  signal VGA_l076_n_220, VGA_l076_n_221, VGA_l076_n_222, VGA_l076_n_223, VGA_l076_n_224 : std_logic;
  signal VGA_l076_n_225, VGA_l076_n_226, VGA_l076_n_227, VGA_l076_n_228, VGA_l076_n_229 : std_logic;
  signal VGA_l076_n_230, VGA_l076_n_231, VGA_l076_n_233, VGA_l076_n_235, VGA_l076_n_236 : std_logic;
  signal VGA_l076_n_237, VGA_l076_n_238, VGA_l076_n_239, VGA_l076_n_241, VGA_l076_n_242 : std_logic;
  signal VGA_l076_n_243, VGA_l0410_n_0, VGA_l0410_n_1, VGA_l0410_n_2, VGA_l0410_n_3 : std_logic;
  signal VGA_l0410_n_4, VGA_l0410_n_5, VGA_l0410_n_6, VGA_l0410_n_7, VGA_l0410_n_8 : std_logic;
  signal VGA_l0410_n_9, VGA_l0410_n_10, VGA_l0410_n_11, VGA_l0410_n_12, VGA_n_0 : std_logic;
  signal VGA_n_1, VGA_n_2, VGA_n_3, VGA_n_4, VGA_n_5 : std_logic;
  signal VGA_n_6, VGA_n_7, VGA_n_8, VGA_r1, VGA_r2 : std_logic;
  signal VGA_r3, VGA_r4, VGA_r5, VGA_r6, VGA_r7 : std_logic;
  signal VGA_r8, VGA_r9, VGA_r10, e_1, e_2 : std_logic;
  signal e_3, e_4, e_5, e_6, n_0 : std_logic;
  signal n_1, n_2, n_3, n_4, n_5 : std_logic;
  signal spawn_or_not_e1, spawn_or_not_e2, spawn_or_not_e3, spawn_or_not_e4, spawn_or_not_e5 : std_logic;
  signal spawn_or_not_e6 : std_logic;

begin

  Movement_module : movement port map(clk => clk, reset => reset, frame_ready => n_5, left => left, right => right, up => up, down => down, shoot => shoot, enemy_1_y(8) => y_e_spawn_1(8:7), enemy_1_y(7) => n_4, enemy_1_y(6) => y_e_spawn_1(5:0), enemy_2_y(8) => y_e_spawn_1(8), enemy_2_y(7) => y_e_spawn_2(7), enemy_2_y(6) => n_4, enemy_2_y(5) => y_e_spawn_1(7), enemy_2_y(4) => y_e_spawn_1(4), enemy_2_y(3) => y_e_spawn_2(3), enemy_2_y(2) => y_e_spawn_1(3), enemy_2_y(1) => y_e_spawn_2(1), enemy_2_y(0) => y_e_spawn_2(1), enemy_3_y(8) => y_e_spawn_1(5), enemy_3_y(7) => y_e_spawn_3(7), enemy_3_y(6) => n_2, enemy_3_y(5) => y_e_spawn_1(4), enemy_3_y(4) => y_e_spawn_1(2), enemy_3_y(3) => y_e_spawn_3(3), enemy_3_y(2) => y_e_spawn_1(1), enemy_3_y(1) => y_e_spawn_3(1), enemy_3_y(0) => y_e_spawn_1(0), enemy_4_y(8) => y_e_spawn_2(7), enemy_4_y(7) => y_e_spawn_4(7), enemy_4_y(6) => n_0, enemy_4_y(5) => y_e_spawn_1(5:4), enemy_4_y(4) => y_e_spawn_2(1), enemy_4_y(3) => y_e_spawn_1(2), enemy_4_y(2) => y_e_spawn_3(1), enemy_4_y(1) => y_e_spawn_1(1), enemy_5_y(8) => y_e_spawn_5(8), enemy_5_y(7) => y_e_spawn_2(7), enemy_5_y(6) => n_1, enemy_5_y(5) => y_e_spawn_1(7), enemy_5_y(4) => y_e_spawn_1(5), enemy_5_y(3) => y_e_spawn_1(3), enemy_5_y(2) => y_e_spawn_3(3), enemy_5_y(1) => y_e_spawn_1(1), enemy_5_y(0) => y_e_spawn_2(1), enemy_6_y(8) => y_e_spawn_2(1), enemy_6_y(7) => y_e_spawn_3(1), enemy_6_y(6) => n_3, enemy_6_y(5) => y_e_spawn_1(1), enemy_6_y(4) => y_e_spawn_1(4), enemy_6_y(3) => y_e_spawn_3(7), enemy_6_y(2) => y_e_spawn_1(2), enemy_6_y(1) => y_e_spawn_2(7), enemy_6_y(0) => y_e_spawn_5(8), e_respawn_1 => spawn_or_not_e1, e_respawn_2 => spawn_or_not_e2, e_respawn_3 => spawn_or_not_e3, e_respawn_4 => spawn_or_not_e4, e_respawn_5 => spawn_or_not_e5, e_respawn_6 => spawn_or_not_e6, coll_enemy_1 => collision_output_vector(9), coll_enemy_2 => collision_output_vector(10), coll_enemy_3 => collision_output_vector(11), coll_enemy_4 => collision_output_vector(12), coll_enemy_5 => collision_output_vector(13), coll_enemy_6 => collision_output_vector(14), coll_bullet_1 => collision_output_vector(0), coll_bullet_2 => collision_output_vector(1), coll_bullet_3 => collision_output_vector(2), coll_player => collision_output_vector(4), player_x => x_pos_p, player_y => y_pos_p, enemy_x_1 => x_pos_e1, enemy_y_1 => y_pos_e1, enemy_x_2 => x_pos_e2, enemy_y_2 => y_pos_e2, enemy_x_3 => x_pos_e3, enemy_y_3 => y_pos_e3, enemy_x_4 => x_pos_e4, enemy_y_4 => y_pos_e4, enemy_x_5 => x_pos_e5, enemy_y_5 => y_pos_e5, enemy_x_6 => x_pos_e6, enemy_y_6 => y_pos_e6, bullet_x_1 => x_pos_b1, bullet_y_1 => y_pos_b1, bullet_x_2 => x_pos_b2, bullet_y_2 => y_pos_b2, bullet_x_3 => x_pos_b3, bullet_y_3 => y_pos_b3, enemy_alive_1 => e_1, enemy_alive_2 => e_2, enemy_alive_3 => e_3, enemy_alive_4 => e_4, enemy_alive_5 => e_5, enemy_alive_6 => e_6);
  g12 : INVD0BWP7T port map(I => v_sync, ZN => n_5);
  g11 : INVD0BWP7T port map(I => y_e_spawn_2(1), ZN => n_3);
  g8 : INVD0BWP7T port map(I => y_e_spawn_1(5), ZN => n_2);
  g7 : INVD0BWP7T port map(I => y_e_spawn_1(8), ZN => n_4);
  g9 : INVD0BWP7T port map(I => y_e_spawn_5(8), ZN => n_1);
  g10 : INVD0BWP7T port map(I => y_e_spawn_2(7), ZN => n_0);
  VGA_g112 : ND2D4BWP7T port map(A1 => VGA_n_8, A2 => VGA_n_7, ZN => r);
  VGA_g113 : INR3D0BWP7T port map(A1 => VGA_n_6, B1 => VGA_r3, B2 => VGA_r4, ZN => VGA_n_8);
  VGA_g114 : NR4D0BWP7T port map(A1 => VGA_r10, A2 => VGA_r9, A3 => VGA_r6, A4 => VGA_r5, ZN => VGA_n_7);
  VGA_g115 : NR4D0BWP7T port map(A1 => VGA_r8, A2 => VGA_r7, A3 => VGA_r1, A4 => VGA_r2, ZN => VGA_n_6);
  VGA_g116 : ND2D4BWP7T port map(A1 => VGA_n_5, A2 => VGA_n_4, ZN => g);
  VGA_g117 : INR3D0BWP7T port map(A1 => VGA_n_3, B1 => VGA_g3, B2 => VGA_g4, ZN => VGA_n_5);
  VGA_g118 : NR4D0BWP7T port map(A1 => VGA_g5, A2 => VGA_g6, A3 => VGA_g9, A4 => VGA_g10, ZN => VGA_n_4);
  VGA_g119 : NR4D0BWP7T port map(A1 => VGA_g7, A2 => VGA_g8, A3 => VGA_g2, A4 => VGA_g1, ZN => VGA_n_3);
  VGA_g120 : ND2D4BWP7T port map(A1 => VGA_n_2, A2 => VGA_n_1, ZN => b);
  VGA_g121 : INR3D0BWP7T port map(A1 => VGA_n_0, B1 => VGA_b3, B2 => VGA_b4, ZN => VGA_n_2);
  VGA_g122 : NR4D0BWP7T port map(A1 => VGA_b10, A2 => VGA_b9, A3 => VGA_b6, A4 => VGA_b5, ZN => VGA_n_1);
  VGA_g123 : NR4D0BWP7T port map(A1 => VGA_b8, A2 => VGA_b7, A3 => VGA_b2, A4 => VGA_b1, ZN => VGA_n_0);
  VGA_l071_g12402 : OAI211D0BWP7T port map(A1 => VGA_l071_n_76, A2 => VGA_l071_n_195, B => VGA_l071_n_243, C => VGA_l071_n_223, ZN => VGA_r5);
  VGA_l071_g12403 : AOI211D0BWP7T port map(A1 => VGA_l071_n_206, A2 => VGA_l071_n_111, B => VGA_l071_n_242, C => VGA_l071_n_225, ZN => VGA_l071_n_243);
  VGA_l071_g12404 : OAI211D0BWP7T port map(A1 => VGA_l071_n_162, A2 => VGA_l071_n_216, B => VGA_l071_n_241, C => VGA_l071_n_238, ZN => VGA_l071_n_242);
  VGA_l071_g12405 : NR4D0BWP7T port map(A1 => VGA_l071_n_239, A2 => VGA_l071_n_227, A3 => VGA_l071_n_219, A4 => VGA_l071_n_220, ZN => VGA_l071_n_241);
  VGA_l071_g12406 : OAI211D0BWP7T port map(A1 => VGA_l071_n_91, A2 => VGA_l071_n_212, B => VGA_l071_n_237, C => VGA_l071_n_235, ZN => VGA_g5);
  VGA_l071_g12407 : NR4D0BWP7T port map(A1 => VGA_l071_n_233, A2 => VGA_l071_n_191, A3 => VGA_l071_n_151, A4 => VGA_l071_n_138, ZN => VGA_l071_n_239);
  VGA_l071_g12408 : NR4D0BWP7T port map(A1 => VGA_l071_n_226, A2 => VGA_l071_n_228, A3 => VGA_l071_n_221, A4 => VGA_l071_n_192, ZN => VGA_l071_n_238);
  VGA_l071_g12409 : AOI211D0BWP7T port map(A1 => VGA_l071_n_206, A2 => VGA_l071_n_117, B => VGA_l071_n_236, C => VGA_l071_n_218, ZN => VGA_l071_n_237);
  VGA_l071_g12410 : OAI211D0BWP7T port map(A1 => VGA_l071_n_99, A2 => VGA_l071_n_195, B => VGA_l071_n_230, C => VGA_l071_n_224, ZN => VGA_l071_n_236);
  VGA_l071_g12411 : AOI211D0BWP7T port map(A1 => VGA_l071_n_211, A2 => VGA_l071_n_137, B => VGA_l071_n_231, C => VGA_l071_n_213, ZN => VGA_l071_n_235);
  VGA_l071_g12412 : OAI32D0BWP7T port map(A1 => VGA_l071_n_24, A2 => VGA_l071_n_60, A3 => VGA_l071_n_216, B1 => VGA_l071_n_94, B2 => VGA_l071_n_215, ZN => VGA_b5);
  VGA_l071_g12413 : ND4D0BWP7T port map(A1 => VGA_l071_n_210, A2 => VGA_l071_n_189, A3 => VGA_l071_n_176, A4 => VGA_l071_n_165, ZN => VGA_l071_n_233);
  VGA_l071_g12414 : OAI211D0BWP7T port map(A1 => VGA_l071_n_191, A2 => VGA_l071_n_209, B => VGA_l071_n_204, C => VGA_l071_n_199, ZN => VGA_enable5);
  VGA_l071_g12415 : OAI22D0BWP7T port map(A1 => VGA_l071_n_217, A2 => VGA_l071_n_139, B1 => VGA_l071_n_207, B2 => VGA_l071_n_131, ZN => VGA_l071_n_231);
  VGA_l071_g12416 : AOI31D0BWP7T port map(A1 => VGA_l071_n_190, A2 => VGA_l071_n_182, A3 => VGA_l071_n_77, B => VGA_l071_n_229, ZN => VGA_l071_n_230);
  VGA_l071_g12417 : AOI21D0BWP7T port map(A1 => VGA_l071_n_103, A2 => VGA_l071_n_86, B => VGA_l071_n_216, ZN => VGA_l071_n_229);
  VGA_l071_g12418 : AOI31D0BWP7T port map(A1 => VGA_l071_n_145, A2 => VGA_l071_n_88, A3 => VGA_l071_n_75, B => VGA_l071_n_217, ZN => VGA_l071_n_228);
  VGA_l071_g12419 : AOI31D0BWP7T port map(A1 => VGA_l071_n_122, A2 => VGA_l071_n_118, A3 => VGA_l071_n_60, B => VGA_l071_n_214, ZN => VGA_l071_n_227);
  VGA_l071_g12420 : AOI31D0BWP7T port map(A1 => VGA_l071_n_142, A2 => VGA_l071_n_122, A3 => VGA_l071_n_88, B => VGA_l071_n_215, ZN => VGA_l071_n_226);
  VGA_l071_g12421 : AOI22D0BWP7T port map(A1 => VGA_l071_n_205, A2 => VGA_l071_n_195, B1 => VGA_l071_n_119, B2 => VGA_l071_n_89, ZN => VGA_l071_n_225);
  VGA_l071_g12422 : AO21D0BWP7T port map(A1 => VGA_l071_n_123, A2 => VGA_l071_n_91, B => VGA_l071_n_215, Z => VGA_l071_n_224);
  VGA_l071_g12423 : OA21D0BWP7T port map(A1 => VGA_l071_n_208, A2 => VGA_l071_n_157, B => VGA_l071_n_222, Z => VGA_l071_n_223);
  VGA_l071_g12424 : AO31D0BWP7T port map(A1 => VGA_l071_n_135, A2 => VGA_l071_n_68, A3 => VGA_l071_n_69, B => VGA_l071_n_204, Z => VGA_l071_n_222);
  VGA_l071_g12425 : AOI21D0BWP7T port map(A1 => VGA_l071_n_89, A2 => VGA_l071_n_52, B => VGA_l071_n_212, ZN => VGA_l071_n_221);
  VGA_l071_g12426 : AOI31D0BWP7T port map(A1 => VGA_l071_n_132, A2 => VGA_l071_n_76, A3 => VGA_l071_n_58, B => VGA_l071_n_207, ZN => VGA_l071_n_220);
  VGA_l071_g12427 : OA21D0BWP7T port map(A1 => VGA_l071_n_134, A2 => VGA_l071_n_90, B => VGA_l071_n_211, Z => VGA_l071_n_219);
  VGA_l071_g12428 : AOI21D0BWP7T port map(A1 => VGA_l071_n_88, A2 => VGA_l071_n_0, B => VGA_l071_n_204, ZN => VGA_l071_n_218);
  VGA_l071_g12429 : AOI32D0BWP7T port map(A1 => VGA_l071_n_190, A2 => VGA_l071_n_181, A3 => VGA_l071_n_38, B1 => VGA_l071_n_202, B2 => VGA_l071_n_154, ZN => VGA_l071_n_214);
  VGA_l071_g12430 : AOI21D0BWP7T port map(A1 => VGA_l071_n_103, A2 => VGA_l071_n_68, B => VGA_l071_n_208, ZN => VGA_l071_n_213);
  VGA_l071_g12431 : AOI22D0BWP7T port map(A1 => VGA_l071_n_203, A2 => VGA_l071_n_156, B1 => VGA_l071_n_202, B2 => VGA_l071_n_143, ZN => VGA_l071_n_217);
  VGA_l071_g12432 : AOI22D0BWP7T port map(A1 => VGA_l071_n_202, A2 => VGA_l071_n_160, B1 => VGA_l071_n_203, B2 => VGA_l071_n_144, ZN => VGA_l071_n_216);
  VGA_l071_g12433 : AOI32D0BWP7T port map(A1 => VGA_l071_n_198, A2 => VGA_l071_n_1, A3 => VGA_l071_n_104, B1 => VGA_l071_n_203, B2 => VGA_l071_n_155, ZN => VGA_l071_n_215);
  VGA_l071_g12434 : OAI31D0BWP7T port map(A1 => VGA_l071_n_2, A2 => VGA_l071_n_127, A3 => VGA_l071_n_179, B => VGA_l071_n_201, ZN => VGA_l071_n_210);
  VGA_l071_g12435 : NR4D0BWP7T port map(A1 => VGA_l071_n_200, A2 => VGA_l071_n_186, A3 => VGA_l071_n_182, A4 => VGA_l071_n_185, ZN => VGA_l071_n_209);
  VGA_l071_g12436 : MAOI22D0BWP7T port map(A1 => VGA_l071_n_196, A2 => VGA_l071_n_170, B1 => VGA_l071_n_191, B2 => VGA_l071_n_165, ZN => VGA_l071_n_212);
  VGA_l071_g12437 : OAI22D0BWP7T port map(A1 => VGA_l071_n_197, A2 => VGA_l071_n_171, B1 => VGA_l071_n_193, B2 => VGA_l071_n_150, ZN => VGA_l071_n_211);
  VGA_l071_g12438 : CKND1BWP7T port map(I => VGA_l071_n_206, ZN => VGA_l071_n_205);
  VGA_l071_g12439 : AOI22D0BWP7T port map(A1 => VGA_l071_n_196, A2 => VGA_l071_n_169, B1 => VGA_l071_n_194, B2 => VGA_l071_n_151, ZN => VGA_l071_n_208);
  VGA_l071_g12440 : MAOI22D0BWP7T port map(A1 => VGA_l071_n_196, A2 => VGA_l071_n_151, B1 => VGA_l071_n_193, B2 => VGA_l071_n_168, ZN => VGA_l071_n_207);
  VGA_l071_g12441 : OAI22D0BWP7T port map(A1 => VGA_l071_n_197, A2 => VGA_l071_n_167, B1 => VGA_l071_n_191, B2 => VGA_l071_n_176, ZN => VGA_l071_n_206);
  VGA_l071_g12442 : MAOI22D0BWP7T port map(A1 => VGA_l071_n_196, A2 => VGA_l071_n_140, B1 => VGA_l071_n_193, B2 => VGA_l071_n_167, ZN => VGA_l071_n_204);
  VGA_l071_g12443 : INR2D0BWP7T port map(A1 => VGA_l071_n_198, B1 => VGA_l071_n_114, ZN => VGA_l071_n_203);
  VGA_l071_g12444 : INR2D0BWP7T port map(A1 => VGA_l071_n_198, B1 => VGA_l071_n_113, ZN => VGA_l071_n_202);
  VGA_l071_g12445 : CKND1BWP7T port map(I => VGA_l071_n_200, ZN => VGA_l071_n_201);
  VGA_l071_g12446 : OAI21D0BWP7T port map(A1 => VGA_l071_n_177, A2 => VGA_l071_n_161, B => VGA_l071_n_194, ZN => VGA_l071_n_199);
  VGA_l071_g12447 : ND3D0BWP7T port map(A1 => VGA_l071_n_188, A2 => VGA_l071_n_176, A3 => VGA_l071_n_165, ZN => VGA_l071_n_200);
  VGA_l071_g12448 : INVD0BWP7T port map(I => VGA_l071_n_197, ZN => VGA_l071_n_196);
  VGA_l071_g12449 : INR2D0BWP7T port map(A1 => VGA_l071_n_185, B1 => VGA_l071_n_191, ZN => VGA_l071_n_198);
  VGA_l071_g12450 : ND2D0BWP7T port map(A1 => VGA_l071_n_190, A2 => VGA_l071_n_184, ZN => VGA_l071_n_197);
  VGA_l071_g12451 : CKND1BWP7T port map(I => VGA_l071_n_193, ZN => VGA_l071_n_194);
  VGA_l071_g12452 : AOI211D0BWP7T port map(A1 => VGA_l071_n_122, A2 => VGA_l071_n_74, B => VGA_l071_n_191, C => VGA_l071_n_183, ZN => VGA_l071_n_192);
  VGA_l071_g12453 : IND2D0BWP7T port map(A1 => VGA_l071_n_189, B1 => VGA_l071_n_190, ZN => VGA_l071_n_195);
  VGA_l071_g12454 : ND2D0BWP7T port map(A1 => VGA_l071_n_190, A2 => VGA_l071_n_164, ZN => VGA_l071_n_193);
  VGA_l071_g12455 : INVD1BWP7T port map(I => VGA_l071_n_191, ZN => VGA_l071_n_190);
  VGA_l071_g12456 : OAI221D0BWP7T port map(A1 => VGA_l071_n_49, A2 => VGA_l071_n_32, B1 => VGA_l071_n_20, B2 => VGA_l071_n_21, C => VGA_l071_n_187, ZN => VGA_l071_n_191);
  VGA_l071_g12457 : AOI22D0BWP7T port map(A1 => VGA_l071_n_184, A2 => VGA_l071_n_161, B1 => VGA_l071_n_170, B2 => VGA_l071_n_164, ZN => VGA_l071_n_188);
  VGA_l071_g12458 : AOI33D0BWP7T port map(A1 => VGA_l071_n_184, A2 => VGA_l071_n_143, A3 => VGA_l071_n_113, B1 => VGA_l071_n_164, B2 => VGA_l071_n_156, B3 => VGA_l071_n_114, ZN => VGA_l071_n_189);
  VGA_l071_g12459 : AOI211D0BWP7T port map(A1 => VGA_l071_n_173, A2 => VGA_l071_n_136, B => VGA_l071_n_178, C => VGA_l071_n_120, ZN => VGA_l071_n_187);
  VGA_l071_g12460 : OA21D0BWP7T port map(A1 => VGA_l071_n_180, A2 => VGA_l071_n_170, B => VGA_l071_n_184, Z => VGA_l071_n_186);
  VGA_l071_g12461 : NR2D0BWP7T port map(A1 => VGA_l071_n_179, A2 => VGA_l071_n_115, ZN => VGA_l071_n_185);
  VGA_l071_g12462 : NR2D0BWP7T port map(A1 => VGA_l071_n_179, A2 => VGA_l071_n_116, ZN => VGA_l071_n_184);
  VGA_l071_g12463 : CKND1BWP7T port map(I => VGA_l071_n_182, ZN => VGA_l071_n_183);
  VGA_l071_g12464 : AO32D0BWP7T port map(A1 => VGA_l071_n_166, A2 => VGA_l071_n_102, A3 => VGA_l071_n_37, B1 => VGA_l071_n_175, B2 => VGA_y(4), Z => VGA_l071_n_181);
  VGA_l071_g12465 : OAI22D0BWP7T port map(A1 => VGA_l071_n_172, A2 => VGA_l071_n_113, B1 => VGA_l071_n_174, B2 => VGA_l071_n_38, ZN => VGA_l071_n_182);
  VGA_l071_g12466 : IND2D0BWP7T port map(A1 => VGA_l071_n_177, B1 => VGA_l071_n_167, ZN => VGA_l071_n_180);
  VGA_l071_g12467 : MOAI22D0BWP7T port map(A1 => VGA_l071_n_163, A2 => VGA_l071_n_136, B1 => VGA_l071_n_21, B2 => VGA_l071_n_20, ZN => VGA_l071_n_178);
  VGA_l071_g12468 : AOI22D0BWP7T port map(A1 => VGA_l071_n_166, A2 => y_pos_e1(4), B1 => VGA_l071_n_159, B2 => VGA_l071_n_11, ZN => VGA_l071_n_179);
  VGA_l071_g12469 : ND2D0BWP7T port map(A1 => VGA_l071_n_168, A2 => VGA_l071_n_171, ZN => VGA_l071_n_177);
  VGA_l071_g12470 : ND2D0BWP7T port map(A1 => VGA_l071_n_164, A2 => VGA_l071_n_140, ZN => VGA_l071_n_176);
  VGA_l071_g12471 : CKND1BWP7T port map(I => VGA_l071_n_174, ZN => VGA_l071_n_175);
  VGA_l071_g12472 : OAI211D0BWP7T port map(A1 => VGA_l071_n_96, A2 => VGA_l071_n_129, B => VGA_l071_n_153, C => VGA_l071_n_105, ZN => VGA_l071_n_173);
  VGA_l071_g12473 : ND3D0BWP7T port map(A1 => VGA_l071_n_154, A2 => VGA_l071_n_158, A3 => VGA_l071_n_115, ZN => VGA_l071_n_172);
  VGA_l071_g12474 : ND3D0BWP7T port map(A1 => VGA_l071_n_159, A2 => VGA_l071_n_102, A3 => VGA_l071_n_37, ZN => VGA_l071_n_174);
  VGA_l071_g12475 : CKND1BWP7T port map(I => VGA_l071_n_168, ZN => VGA_l071_n_169);
  VGA_l071_g12476 : ND2D0BWP7T port map(A1 => VGA_l071_n_156, A2 => VGA_l071_n_114, ZN => VGA_l071_n_171);
  VGA_l071_g12477 : AN2D1BWP7T port map(A1 => VGA_l071_n_154, A2 => VGA_l071_n_113, Z => VGA_l071_n_170);
  VGA_l071_g12478 : ND2D0BWP7T port map(A1 => VGA_l071_n_160, A2 => VGA_l071_n_113, ZN => VGA_l071_n_168);
  VGA_l071_g12479 : ND2D0BWP7T port map(A1 => VGA_l071_n_155, A2 => VGA_l071_n_114, ZN => VGA_l071_n_167);
  VGA_l071_g12480 : AOI221D0BWP7T port map(A1 => VGA_l071_n_125, A2 => VGA_l071_n_95, B1 => VGA_l071_n_45, B2 => VGA_l071_n_81, C => VGA_l071_n_152, ZN => VGA_l071_n_163);
  VGA_l071_g12481 : AN4D1BWP7T port map(A1 => VGA_l071_n_141, A2 => VGA_l071_n_103, A3 => VGA_l071_n_89, A4 => VGA_l071_n_0, Z => VGA_l071_n_162);
  VGA_l071_g12482 : NR3D0BWP7T port map(A1 => VGA_l071_n_149, A2 => VGA_l071_n_44, A3 => VGA_y(4), ZN => VGA_l071_n_166);
  VGA_l071_g12483 : IND3D0BWP7T port map(A1 => VGA_l071_n_127, B1 => VGA_l071_n_2, B2 => VGA_l071_n_158, ZN => VGA_l071_n_165);
  VGA_l071_g12484 : AN2D1BWP7T port map(A1 => VGA_l071_n_158, A2 => VGA_l071_n_116, Z => VGA_l071_n_164);
  VGA_l071_g12485 : IINR4D0BWP7T port map(A1 => VGA_l071_n_122, A2 => VGA_l071_n_69, B1 => VGA_l071_n_133, B2 => VGA_l071_n_77, ZN => VGA_l071_n_157);
  VGA_l071_g12486 : IND2D0BWP7T port map(A1 => VGA_l071_n_151, B1 => VGA_l071_n_150, ZN => VGA_l071_n_161);
  VGA_l071_g12487 : NR3D0BWP7T port map(A1 => VGA_l071_n_148, A2 => VGA_l071_n_87, A3 => VGA_l071_n_40, ZN => VGA_l071_n_160);
  VGA_l071_g12488 : INR2D0BWP7T port map(A1 => VGA_l071_n_44, B1 => VGA_l071_n_149, ZN => VGA_l071_n_159);
  VGA_l071_g12489 : AOI211D0BWP7T port map(A1 => VGA_l071_n_44, A2 => VGA_l071_n_34, B => VGA_l071_n_149, C => VGA_l071_n_98, ZN => VGA_l071_n_158);
  VGA_l071_g12490 : AOI22D0BWP7T port map(A1 => VGA_l071_n_146, A2 => VGA_l071_n_126, B1 => VGA_l071_n_45, B2 => VGA_l071_n_26, ZN => VGA_l071_n_153);
  VGA_l071_g12491 : OAI22D0BWP7T port map(A1 => VGA_l071_n_146, A2 => VGA_l071_n_130, B1 => VGA_l071_n_97, B2 => VGA_x(5), ZN => VGA_l071_n_152);
  VGA_l071_g12492 : INR3D0BWP7T port map(A1 => VGA_l071_n_148, B1 => VGA_l071_n_40, B2 => VGA_l071_n_87, ZN => VGA_l071_n_156);
  VGA_l071_g12493 : AN3D0BWP7T port map(A1 => VGA_l071_n_147, A2 => VGA_l071_n_87, A3 => VGA_l071_n_39, Z => VGA_l071_n_155);
  VGA_l071_g12494 : INR3D0BWP7T port map(A1 => VGA_l071_n_87, B1 => VGA_l071_n_40, B2 => VGA_l071_n_147, ZN => VGA_l071_n_154);
  VGA_l071_g12495 : AN2D1BWP7T port map(A1 => VGA_l071_n_144, A2 => VGA_l071_n_114, Z => VGA_l071_n_151);
  VGA_l071_g12496 : ND2D0BWP7T port map(A1 => VGA_l071_n_143, A2 => VGA_l071_n_113, ZN => VGA_l071_n_150);
  VGA_l071_g12497 : IND4D0BWP7T port map(A1 => VGA_l071_n_108, B1 => VGA_l071_n_109, B2 => VGA_l071_n_106, B3 => VGA_l071_n_107, ZN => VGA_l071_n_149);
  VGA_l071_g12498 : AN3D0BWP7T port map(A1 => VGA_l071_n_128, A2 => VGA_l071_n_70, A3 => VGA_l071_n_76, Z => VGA_l071_n_145);
  VGA_l071_g12499 : OAI221D0BWP7T port map(A1 => VGA_l071_n_101, A2 => y_pos_e1(1), B1 => VGA_l071_n_4, B2 => VGA_l071_n_82, C => VGA_l071_n_100, ZN => VGA_l071_n_148);
  VGA_l071_g12500 : OAI211D0BWP7T port map(A1 => y_pos_e1(1), A2 => VGA_l071_n_41, B => VGA_l071_n_121, C => VGA_l071_n_101, ZN => VGA_l071_n_147);
  VGA_l071_g12501 : MAOI222D0BWP7T port map(A => VGA_x(2), B => x_pos_e1(2), C => VGA_l071_n_83, ZN => VGA_l071_n_146);
  VGA_l071_g12502 : AN3D0BWP7T port map(A1 => VGA_l071_n_124, A2 => VGA_l071_n_94, A3 => VGA_l071_n_92, Z => VGA_l071_n_142);
  VGA_l071_g12503 : INR3D0BWP7T port map(A1 => VGA_l071_n_128, B1 => VGA_l071_n_72, B2 => VGA_l071_n_77, ZN => VGA_l071_n_141);
  VGA_l071_g12504 : AOI211D0BWP7T port map(A1 => VGA_l071_n_101, A2 => VGA_l071_n_100, B => VGA_l071_n_39, C => VGA_l071_n_43, ZN => VGA_l071_n_144);
  VGA_l071_g12505 : AN4D1BWP7T port map(A1 => VGA_l071_n_101, A2 => VGA_l071_n_100, A3 => VGA_l071_n_42, A4 => VGA_l071_n_40, Z => VGA_l071_n_143);
  VGA_l071_g12506 : INR2D0BWP7T port map(A1 => VGA_l071_n_122, B1 => VGA_l071_n_72, ZN => VGA_l071_n_139);
  VGA_l071_g12507 : AN2D1BWP7T port map(A1 => VGA_l071_n_112, A2 => VGA_l071_n_52, Z => VGA_l071_n_138);
  VGA_l071_g12508 : ND2D0BWP7T port map(A1 => VGA_l071_n_123, A2 => VGA_l071_n_131, ZN => VGA_l071_n_137);
  VGA_l071_g12509 : INR2D0BWP7T port map(A1 => VGA_l071_n_104, B1 => VGA_l071_n_1, ZN => VGA_l071_n_140);
  VGA_l071_g12510 : OA221D0BWP7T port map(A1 => VGA_l071_n_67, A2 => VGA_draw_count5(1), B1 => VGA_l071_n_24, B2 => VGA_l071_n_54, C => VGA_l071_n_74, Z => VGA_l071_n_135);
  VGA_l071_g12511 : OAI211D0BWP7T port map(A1 => VGA_draw_count5(1), A2 => VGA_l071_n_58, B => VGA_l071_n_84, C => VGA_l071_n_74, ZN => VGA_l071_n_134);
  VGA_l071_g12512 : OAI211D0BWP7T port map(A1 => VGA_l071_n_13, A2 => VGA_l071_n_54, B => VGA_l071_n_85, C => VGA_l071_n_75, ZN => VGA_l071_n_133);
  VGA_l071_g12513 : OA21D0BWP7T port map(A1 => VGA_l071_n_14, A2 => VGA_l071_n_3, B => VGA_l071_n_124, Z => VGA_l071_n_132);
  VGA_l071_g12514 : ND2D0BWP7T port map(A1 => VGA_l071_n_110, A2 => VGA_l071_n_105, ZN => VGA_l071_n_136);
  VGA_l071_g12515 : CKND1BWP7T port map(I => VGA_l071_n_129, ZN => VGA_l071_n_130);
  VGA_l071_g12516 : CKND1BWP7T port map(I => VGA_l071_n_125, ZN => VGA_l071_n_126);
  VGA_l071_g12517 : IND2D0BWP7T port map(A1 => VGA_l071_n_100, B1 => y_pos_e1(1), ZN => VGA_l071_n_121);
  VGA_l071_g12518 : MOAI22D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l071_n_10, B1 => VGA_l071_n_49, B2 => VGA_l071_n_32, ZN => VGA_l071_n_120);
  VGA_l071_g12519 : AOI21D0BWP7T port map(A1 => VGA_l071_n_59, A2 => VGA_l071_n_27, B => VGA_l071_n_93, ZN => VGA_l071_n_119);
  VGA_l071_g12520 : AOI211D0BWP7T port map(A1 => VGA_l071_n_55, A2 => VGA_l071_n_24, B => VGA_l071_n_93, C => VGA_l071_n_78, ZN => VGA_l071_n_118);
  VGA_l071_g12521 : OAI221D0BWP7T port map(A1 => VGA_l071_n_62, A2 => VGA_l071_n_0, B1 => VGA_l071_n_29, B2 => VGA_l071_n_64, C => VGA_l071_n_92, ZN => VGA_l071_n_117);
  VGA_l071_g12522 : OA21D0BWP7T port map(A1 => VGA_l071_n_62, A2 => VGA_l071_n_64, B => VGA_l071_n_92, Z => VGA_l071_n_131);
  VGA_l071_g12523 : AOI22D0BWP7T port map(A1 => VGA_l071_n_66, A2 => VGA_l071_n_31, B1 => VGA_l071_n_47, B2 => VGA_x(2), ZN => VGA_l071_n_129);
  VGA_l071_g12524 : NR3D0BWP7T port map(A1 => VGA_l071_n_80, A2 => VGA_l071_n_73, A3 => VGA_l071_n_61, ZN => VGA_l071_n_128);
  VGA_l071_g12525 : IND2D0BWP7T port map(A1 => VGA_l071_n_37, B1 => VGA_l071_n_102, ZN => VGA_l071_n_127);
  VGA_l071_g12526 : OAI22D0BWP7T port map(A1 => VGA_l071_n_66, A2 => VGA_l071_n_31, B1 => VGA_l071_n_47, B2 => VGA_x(2), ZN => VGA_l071_n_125);
  VGA_l071_g12527 : AN3D0BWP7T port map(A1 => VGA_l071_n_68, A2 => VGA_l071_n_75, A3 => VGA_l071_n_69, Z => VGA_l071_n_124);
  VGA_l071_g12528 : AN2D1BWP7T port map(A1 => VGA_l071_n_88, A2 => VGA_l071_n_68, Z => VGA_l071_n_123);
  VGA_l071_g12529 : AN2D1BWP7T port map(A1 => VGA_l071_n_89, A2 => VGA_l071_n_58, Z => VGA_l071_n_122);
  VGA_l071_g12530 : AOI221D0BWP7T port map(A1 => VGA_l071_n_61, A2 => VGA_draw_count5(0), B1 => VGA_l071_n_56, B2 => VGA_l071_n_25, C => VGA_l071_n_80, ZN => VGA_l071_n_112);
  VGA_l071_g12531 : AO222D0BWP7T port map(A1 => VGA_l071_n_61, A2 => VGA_l071_n_24, B1 => VGA_l071_n_55, B2 => VGA_l071_n_13, C1 => VGA_l071_n_53, C2 => VGA_l071_n_27, Z => VGA_l071_n_111);
  VGA_l071_g12532 : OAI22D0BWP7T port map(A1 => VGA_l071_n_45, A2 => VGA_l071_n_26, B1 => VGA_l071_n_46, B2 => VGA_l071_n_16, ZN => VGA_l071_n_110);
  VGA_l071_g12533 : MAOI22D0BWP7T port map(A1 => VGA_l071_n_50, A2 => VGA_l071_n_35, B1 => VGA_l071_n_50, B2 => VGA_l071_n_35, ZN => VGA_l071_n_109);
  VGA_l071_g12534 : OAI22D0BWP7T port map(A1 => VGA_l071_n_65, A2 => VGA_l071_n_15, B1 => VGA_l071_n_36, B2 => VGA_y(9), ZN => VGA_l071_n_108);
  VGA_l071_g12535 : AOI22D0BWP7T port map(A1 => VGA_l071_n_65, A2 => VGA_l071_n_15, B1 => VGA_l071_n_36, B2 => VGA_y(9), ZN => VGA_l071_n_107);
  VGA_l071_g12536 : MAOI22D0BWP7T port map(A1 => VGA_l071_n_48, A2 => VGA_l071_n_28, B1 => VGA_l071_n_48, B2 => VGA_l071_n_28, ZN => VGA_l071_n_106);
  VGA_l071_g12538 : MAOI22D0BWP7T port map(A1 => VGA_l071_n_38, A2 => VGA_l071_n_19, B1 => VGA_l071_n_38, B2 => VGA_l071_n_19, ZN => VGA_l071_n_116);
  VGA_l071_g12540 : MOAI22D0BWP7T port map(A1 => VGA_l071_n_38, A2 => VGA_l071_n_22, B1 => VGA_l071_n_38, B2 => VGA_l071_n_22, ZN => VGA_l071_n_115);
  VGA_l071_g12541 : MAOI22D0BWP7T port map(A1 => VGA_l071_n_37, A2 => VGA_l071_n_33, B1 => VGA_l071_n_37, B2 => VGA_l071_n_33, ZN => VGA_l071_n_114);
  VGA_l071_g12542 : MOAI22D0BWP7T port map(A1 => VGA_l071_n_37, A2 => VGA_l071_n_23, B1 => VGA_l071_n_37, B2 => VGA_l071_n_23, ZN => VGA_l071_n_113);
  VGA_l071_g12543 : AOI21D0BWP7T port map(A1 => VGA_l071_n_56, A2 => VGA_l071_n_24, B => VGA_l071_n_63, ZN => VGA_l071_n_99);
  VGA_l071_g12544 : NR2D0BWP7T port map(A1 => VGA_l071_n_44, A2 => VGA_l071_n_34, ZN => VGA_l071_n_98);
  VGA_l071_g12545 : IND2D0BWP7T port map(A1 => VGA_l071_n_46, B1 => x_pos_e1(5), ZN => VGA_l071_n_97);
  VGA_l071_g12546 : ND2D0BWP7T port map(A1 => VGA_l071_n_46, A2 => VGA_l071_n_16, ZN => VGA_l071_n_105);
  VGA_l071_g12547 : NR2D0BWP7T port map(A1 => VGA_l071_n_66, A2 => VGA_l071_n_31, ZN => VGA_l071_n_96);
  VGA_l071_g12548 : NR2D0BWP7T port map(A1 => VGA_l071_n_71, A2 => VGA_l071_n_41, ZN => VGA_l071_n_104);
  VGA_l071_g12550 : NR2D0BWP7T port map(A1 => VGA_l071_n_79, A2 => VGA_l071_n_78, ZN => VGA_l071_n_103);
  VGA_l071_g12551 : NR2D0BWP7T port map(A1 => VGA_l071_n_71, A2 => VGA_l071_n_82, ZN => VGA_l071_n_102);
  VGA_l071_g12552 : ND2D0BWP7T port map(A1 => VGA_l071_n_82, A2 => VGA_y(1), ZN => VGA_l071_n_101);
  VGA_l071_g12553 : IND2D0BWP7T port map(A1 => VGA_y(1), B1 => VGA_l071_n_41, ZN => VGA_l071_n_100);
  VGA_l071_g12554 : CKND1BWP7T port map(I => VGA_l071_n_90, ZN => VGA_l071_n_91);
  VGA_l071_g12555 : AOI21D0BWP7T port map(A1 => VGA_l071_n_59, A2 => VGA_l071_n_25, B => VGA_l071_n_73, ZN => VGA_l071_n_86);
  VGA_l071_g12556 : OAI21D0BWP7T port map(A1 => VGA_l071_n_56, A2 => VGA_l071_n_53, B => VGA_l071_n_24, ZN => VGA_l071_n_85);
  VGA_l071_g12557 : AO21D0BWP7T port map(A1 => VGA_l071_n_60, A2 => VGA_l071_n_54, B => VGA_l071_n_62, Z => VGA_l071_n_84);
  VGA_l071_g12558 : IAO21D0BWP7T port map(A1 => VGA_l071_n_60, A2 => VGA_l071_n_13, B => VGA_l071_n_55, ZN => VGA_l071_n_94);
  VGA_l071_g12559 : OAI21D0BWP7T port map(A1 => VGA_l071_n_52, A2 => VGA_draw_count5(1), B => VGA_l071_n_70, ZN => VGA_l071_n_93);
  VGA_l071_g12560 : AOI22D0BWP7T port map(A1 => VGA_l071_n_51, A2 => VGA_x(0), B1 => VGA_x(1), B2 => VGA_l071_n_6, ZN => VGA_l071_n_83);
  VGA_l071_g12561 : OA22D0BWP7T port map(A1 => VGA_l071_n_64, A2 => VGA_l071_n_12, B1 => VGA_l071_n_25, B2 => VGA_l071_n_0, Z => VGA_l071_n_92);
  VGA_l071_g12562 : OAI21D0BWP7T port map(A1 => VGA_l071_n_57, A2 => VGA_l071_n_13, B => VGA_l071_n_69, ZN => VGA_l071_n_90);
  VGA_l071_g12563 : AOI22D0BWP7T port map(A1 => VGA_l071_n_56, A2 => VGA_l071_n_13, B1 => VGA_l071_n_59, B2 => VGA_l071_n_24, ZN => VGA_l071_n_89);
  VGA_l071_g12564 : IAO21D0BWP7T port map(A1 => VGA_l071_n_0, A2 => VGA_l071_n_24, B => VGA_l071_n_79, ZN => VGA_l071_n_88);
  VGA_l071_g12565 : MOAI22D0BWP7T port map(A1 => VGA_l071_n_43, A2 => VGA_y(0), B1 => VGA_l071_n_43, B2 => VGA_y(0), ZN => VGA_l071_n_87);
  VGA_l071_g12568 : INVD0BWP7T port map(I => VGA_l071_n_41, ZN => VGA_l071_n_82);
  VGA_l071_g12569 : CKND1BWP7T port map(I => VGA_l071_n_26, ZN => VGA_l071_n_81);
  VGA_l071_g12570 : NR2D0BWP7T port map(A1 => VGA_l071_n_54, A2 => VGA_draw_count5(1), ZN => VGA_l071_n_80);
  VGA_l071_g12571 : INR2D0BWP7T port map(A1 => VGA_l071_n_63, B1 => VGA_l071_n_25, ZN => VGA_l071_n_79);
  VGA_l071_g12572 : NR2D0BWP7T port map(A1 => VGA_l071_n_0, A2 => VGA_draw_count5(1), ZN => VGA_l071_n_78);
  VGA_l071_g12573 : NR2D0BWP7T port map(A1 => VGA_l071_n_57, A2 => VGA_l071_n_29, ZN => VGA_l071_n_77);
  VGA_l071_g12574 : ND2D0BWP7T port map(A1 => VGA_l071_n_55, A2 => VGA_draw_count5(1), ZN => VGA_l071_n_76);
  VGA_l071_g12575 : ND2D0BWP7T port map(A1 => VGA_l071_n_53, A2 => VGA_l071_n_13, ZN => VGA_l071_n_75);
  VGA_l071_g12576 : ND2D0BWP7T port map(A1 => VGA_l071_n_53, A2 => VGA_draw_count5(1), ZN => VGA_l071_n_74);
  VGA_l071_g12577 : NR2D0BWP7T port map(A1 => VGA_l071_n_56, A2 => VGA_l071_n_59, ZN => VGA_l071_n_67);
  VGA_l071_g12578 : AN2D1BWP7T port map(A1 => VGA_l071_n_63, A2 => VGA_l071_n_27, Z => VGA_l071_n_73);
  VGA_l071_g12579 : NR2D0BWP7T port map(A1 => VGA_l071_n_52, A2 => VGA_l071_n_13, ZN => VGA_l071_n_72);
  VGA_l071_g12580 : ND2D0BWP7T port map(A1 => VGA_l071_n_40, A2 => VGA_l071_n_43, ZN => VGA_l071_n_71);
  VGA_l071_g12581 : IND2D0BWP7T port map(A1 => VGA_l071_n_62, B1 => VGA_l071_n_56, ZN => VGA_l071_n_70);
  VGA_l071_g12582 : ND2D0BWP7T port map(A1 => VGA_l071_n_63, A2 => VGA_l071_n_13, ZN => VGA_l071_n_69);
  VGA_l071_g12583 : IND2D0BWP7T port map(A1 => VGA_l071_n_62, B1 => VGA_l071_n_63, ZN => VGA_l071_n_68);
  VGA_l071_g12584 : INVD0BWP7T port map(I => VGA_l071_n_61, ZN => VGA_l071_n_60);
  VGA_l071_g12585 : INVD0BWP7T port map(I => VGA_l071_n_59, ZN => VGA_l071_n_58);
  VGA_l071_g12586 : INVD1BWP7T port map(I => VGA_l071_n_57, ZN => VGA_l071_n_56);
  VGA_l071_g12587 : INVD0BWP7T port map(I => VGA_l071_n_55, ZN => VGA_l071_n_54);
  VGA_l071_g12588 : INVD0BWP7T port map(I => VGA_l071_n_53, ZN => VGA_l071_n_52);
  VGA_l071_g12589 : IAO21D0BWP7T port map(A1 => VGA_x(1), A2 => VGA_l071_n_6, B => x_pos_e1(0), ZN => VGA_l071_n_51);
  VGA_l071_g12590 : OAI21D0BWP7T port map(A1 => VGA_l071_n_7, A2 => x_pos_e1(4), B => VGA_l071_n_26, ZN => VGA_l071_n_66);
  VGA_l071_g12591 : AOI21D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l071_n_5, B => VGA_l071_n_28, ZN => VGA_l071_n_65);
  VGA_l071_g12592 : IND2D0BWP7T port map(A1 => VGA_l071_n_30, B1 => VGA_draw_count5(4), ZN => VGA_l071_n_64);
  VGA_l071_g12593 : INR2D0BWP7T port map(A1 => VGA_draw_count5(4), B1 => VGA_l071_n_17, ZN => VGA_l071_n_63);
  VGA_l071_g12594 : INR2D0BWP7T port map(A1 => VGA_l071_n_29, B1 => VGA_l071_n_27, ZN => VGA_l071_n_62);
  VGA_l071_g12596 : NR2D0BWP7T port map(A1 => VGA_l071_n_14, A2 => VGA_draw_count5(4), ZN => VGA_l071_n_61);
  VGA_l071_g12597 : NR2D0BWP7T port map(A1 => VGA_l071_n_30, A2 => VGA_draw_count5(4), ZN => VGA_l071_n_59);
  VGA_l071_g12598 : IND2D0BWP7T port map(A1 => VGA_l071_n_14, B1 => VGA_draw_count5(4), ZN => VGA_l071_n_57);
  VGA_l071_g12599 : NR2D0BWP7T port map(A1 => VGA_l071_n_17, A2 => VGA_draw_count5(4), ZN => VGA_l071_n_55);
  VGA_l071_g12600 : NR2D0BWP7T port map(A1 => VGA_l071_n_18, A2 => VGA_draw_count5(4), ZN => VGA_l071_n_53);
  VGA_l071_g12601 : CKND1BWP7T port map(I => VGA_l071_n_43, ZN => VGA_l071_n_42);
  VGA_l071_g12602 : CKND1BWP7T port map(I => VGA_l071_n_40, ZN => VGA_l071_n_39);
  VGA_l071_g12603 : MOAI22D0BWP7T port map(A1 => VGA_y(8), A2 => y_pos_e1(8), B1 => VGA_y(8), B2 => y_pos_e1(8), ZN => VGA_l071_n_50);
  VGA_l071_g12604 : MOAI22D0BWP7T port map(A1 => VGA_x(7), A2 => x_pos_e1(7), B1 => VGA_x(7), B2 => x_pos_e1(7), ZN => VGA_l071_n_49);
  VGA_l071_g12605 : MOAI22D0BWP7T port map(A1 => VGA_y(7), A2 => y_pos_e1(7), B1 => VGA_y(7), B2 => y_pos_e1(7), ZN => VGA_l071_n_48);
  VGA_l071_g12606 : MAOI22D0BWP7T port map(A1 => VGA_x(3), A2 => x_pos_e1(3), B1 => VGA_x(3), B2 => x_pos_e1(3), ZN => VGA_l071_n_47);
  VGA_l071_g12607 : MOAI22D0BWP7T port map(A1 => VGA_x(6), A2 => x_pos_e1(6), B1 => VGA_x(6), B2 => x_pos_e1(6), ZN => VGA_l071_n_46);
  VGA_l071_g12608 : MOAI22D0BWP7T port map(A1 => VGA_x(5), A2 => x_pos_e1(5), B1 => VGA_x(5), B2 => x_pos_e1(5), ZN => VGA_l071_n_45);
  VGA_l071_g12609 : MAOI22D0BWP7T port map(A1 => VGA_y(5), A2 => y_pos_e1(5), B1 => VGA_y(5), B2 => y_pos_e1(5), ZN => VGA_l071_n_44);
  VGA_l071_g12610 : MOAI22D0BWP7T port map(A1 => VGA_y(1), A2 => y_pos_e1(1), B1 => VGA_y(1), B2 => y_pos_e1(1), ZN => VGA_l071_n_43);
  VGA_l071_g12611 : MOAI22D0BWP7T port map(A1 => VGA_y(2), A2 => y_pos_e1(2), B1 => VGA_y(2), B2 => y_pos_e1(2), ZN => VGA_l071_n_41);
  VGA_l071_g12612 : MOAI22D0BWP7T port map(A1 => VGA_y(0), A2 => y_pos_e1(0), B1 => VGA_y(0), B2 => y_pos_e1(0), ZN => VGA_l071_n_40);
  VGA_l071_g12613 : MAOI22D0BWP7T port map(A1 => VGA_y(4), A2 => y_pos_e1(4), B1 => VGA_y(4), B2 => y_pos_e1(4), ZN => VGA_l071_n_38);
  VGA_l071_g12614 : MOAI22D0BWP7T port map(A1 => VGA_y(3), A2 => y_pos_e1(3), B1 => VGA_y(3), B2 => y_pos_e1(3), ZN => VGA_l071_n_37);
  VGA_l071_g12615 : INVD1BWP7T port map(I => VGA_l071_n_25, ZN => VGA_l071_n_24);
  VGA_l071_g12616 : IND2D0BWP7T port map(A1 => VGA_y(8), B1 => y_pos_e1(8), ZN => VGA_l071_n_36);
  VGA_l071_g12617 : INR2D0BWP7T port map(A1 => y_pos_e1(7), B1 => VGA_y(7), ZN => VGA_l071_n_35);
  VGA_l071_g12618 : IND2D0BWP7T port map(A1 => y_pos_e1(4), B1 => VGA_y(4), ZN => VGA_l071_n_34);
  VGA_l071_g12619 : IND2D0BWP7T port map(A1 => y_pos_e1(2), B1 => VGA_y(2), ZN => VGA_l071_n_33);
  VGA_l071_g12620 : IND2D0BWP7T port map(A1 => x_pos_e1(6), B1 => VGA_x(6), ZN => VGA_l071_n_32);
  VGA_l071_g12621 : IND2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_e1(3), ZN => VGA_l071_n_31);
  VGA_l071_g12622 : ND2D0BWP7T port map(A1 => VGA_draw_count5(2), A2 => VGA_draw_count5(3), ZN => VGA_l071_n_30);
  VGA_l071_g12623 : ND2D0BWP7T port map(A1 => VGA_l071_n_3, A2 => VGA_draw_count5(0), ZN => VGA_l071_n_29);
  VGA_l071_g12624 : NR2D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l071_n_5, ZN => VGA_l071_n_28);
  VGA_l071_g12625 : NR2D0BWP7T port map(A1 => VGA_l071_n_3, A2 => VGA_draw_count5(0), ZN => VGA_l071_n_27);
  VGA_l071_g12626 : ND2D0BWP7T port map(A1 => VGA_l071_n_7, A2 => x_pos_e1(4), ZN => VGA_l071_n_26);
  VGA_l071_g12627 : ND2D0BWP7T port map(A1 => VGA_draw_count5(1), A2 => VGA_draw_count5(0), ZN => VGA_l071_n_25);
  VGA_l071_g12629 : CKND1BWP7T port map(I => VGA_l071_n_13, ZN => VGA_l071_n_12);
  VGA_l071_g12630 : IND2D0BWP7T port map(A1 => VGA_y(4), B1 => y_pos_e1(4), ZN => VGA_l071_n_11);
  VGA_l071_g12631 : ND2D0BWP7T port map(A1 => VGA_l071_n_8, A2 => y_pos_e1(2), ZN => VGA_l071_n_23);
  VGA_l071_g12632 : NR2D0BWP7T port map(A1 => VGA_l071_n_9, A2 => y_pos_e1(3), ZN => VGA_l071_n_22);
  VGA_l071_g12633 : INR2D0BWP7T port map(A1 => x_pos_e1(7), B1 => VGA_x(7), ZN => VGA_l071_n_21);
  VGA_l071_g12634 : ND2D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l071_n_10, ZN => VGA_l071_n_20);
  VGA_l071_g12635 : INR2D0BWP7T port map(A1 => y_pos_e1(3), B1 => VGA_y(3), ZN => VGA_l071_n_19);
  VGA_l071_g12636 : IND2D0BWP7T port map(A1 => VGA_draw_count5(2), B1 => VGA_draw_count5(3), ZN => VGA_l071_n_18);
  VGA_l071_g12637 : IND2D0BWP7T port map(A1 => VGA_draw_count5(3), B1 => VGA_draw_count5(2), ZN => VGA_l071_n_17);
  VGA_l071_g12638 : INR2D0BWP7T port map(A1 => VGA_x(5), B1 => x_pos_e1(5), ZN => VGA_l071_n_16);
  VGA_l071_g12639 : IND2D0BWP7T port map(A1 => y_pos_e1(5), B1 => VGA_y(5), ZN => VGA_l071_n_15);
  VGA_l071_g12640 : OR2D0BWP7T port map(A1 => VGA_draw_count5(2), A2 => VGA_draw_count5(3), Z => VGA_l071_n_14);
  VGA_l071_g12641 : NR2D0BWP7T port map(A1 => VGA_draw_count5(1), A2 => VGA_draw_count5(0), ZN => VGA_l071_n_13);
  VGA_l071_g12642 : CKND1BWP7T port map(I => x_pos_e1(8), ZN => VGA_l071_n_10);
  VGA_l071_g12643 : CKND1BWP7T port map(I => VGA_y(3), ZN => VGA_l071_n_9);
  VGA_l071_g12644 : CKND1BWP7T port map(I => VGA_y(2), ZN => VGA_l071_n_8);
  VGA_l071_g12645 : CKND1BWP7T port map(I => VGA_x(4), ZN => VGA_l071_n_7);
  VGA_l071_g12646 : CKND1BWP7T port map(I => x_pos_e1(1), ZN => VGA_l071_n_6);
  VGA_l071_g12647 : CKND1BWP7T port map(I => y_pos_e1(6), ZN => VGA_l071_n_5);
  VGA_l071_g12648 : CKND1BWP7T port map(I => y_pos_e1(1), ZN => VGA_l071_n_4);
  VGA_l071_g12649 : INVD0BWP7T port map(I => VGA_draw_count5(1), ZN => VGA_l071_n_3);
  VGA_l071_g2 : MUX2ND0BWP7T port map(I0 => VGA_y(3), I1 => VGA_l071_n_9, S => VGA_l071_n_38, ZN => VGA_l071_n_2);
  VGA_l071_g12650 : MUX2ND0BWP7T port map(I0 => VGA_l071_n_8, I1 => VGA_y(2), S => VGA_l071_n_37, ZN => VGA_l071_n_1);
  VGA_l071_g12651 : IND2D1BWP7T port map(A1 => VGA_l071_n_18, B1 => VGA_draw_count5(4), ZN => VGA_l071_n_0);
  VGA_l071_g12652 : INVD0BWP7T port map(I => VGA_l071_n_66, ZN => VGA_l071_n_95);
  VGA_l072_g12402 : OAI211D0BWP7T port map(A1 => VGA_l072_n_76, A2 => VGA_l072_n_195, B => VGA_l072_n_243, C => VGA_l072_n_223, ZN => VGA_r6);
  VGA_l072_g12403 : AOI211D0BWP7T port map(A1 => VGA_l072_n_206, A2 => VGA_l072_n_111, B => VGA_l072_n_242, C => VGA_l072_n_225, ZN => VGA_l072_n_243);
  VGA_l072_g12404 : OAI211D0BWP7T port map(A1 => VGA_l072_n_162, A2 => VGA_l072_n_216, B => VGA_l072_n_241, C => VGA_l072_n_238, ZN => VGA_l072_n_242);
  VGA_l072_g12405 : NR4D0BWP7T port map(A1 => VGA_l072_n_239, A2 => VGA_l072_n_227, A3 => VGA_l072_n_219, A4 => VGA_l072_n_220, ZN => VGA_l072_n_241);
  VGA_l072_g12406 : OAI211D0BWP7T port map(A1 => VGA_l072_n_91, A2 => VGA_l072_n_212, B => VGA_l072_n_237, C => VGA_l072_n_235, ZN => VGA_g6);
  VGA_l072_g12407 : NR4D0BWP7T port map(A1 => VGA_l072_n_233, A2 => VGA_l072_n_191, A3 => VGA_l072_n_151, A4 => VGA_l072_n_138, ZN => VGA_l072_n_239);
  VGA_l072_g12408 : NR4D0BWP7T port map(A1 => VGA_l072_n_226, A2 => VGA_l072_n_228, A3 => VGA_l072_n_221, A4 => VGA_l072_n_192, ZN => VGA_l072_n_238);
  VGA_l072_g12409 : AOI211D0BWP7T port map(A1 => VGA_l072_n_206, A2 => VGA_l072_n_117, B => VGA_l072_n_236, C => VGA_l072_n_218, ZN => VGA_l072_n_237);
  VGA_l072_g12410 : OAI211D0BWP7T port map(A1 => VGA_l072_n_99, A2 => VGA_l072_n_195, B => VGA_l072_n_230, C => VGA_l072_n_224, ZN => VGA_l072_n_236);
  VGA_l072_g12411 : AOI211D0BWP7T port map(A1 => VGA_l072_n_211, A2 => VGA_l072_n_137, B => VGA_l072_n_231, C => VGA_l072_n_213, ZN => VGA_l072_n_235);
  VGA_l072_g12412 : OAI32D0BWP7T port map(A1 => VGA_l072_n_24, A2 => VGA_l072_n_60, A3 => VGA_l072_n_216, B1 => VGA_l072_n_94, B2 => VGA_l072_n_215, ZN => VGA_b6);
  VGA_l072_g12413 : ND4D0BWP7T port map(A1 => VGA_l072_n_210, A2 => VGA_l072_n_189, A3 => VGA_l072_n_176, A4 => VGA_l072_n_165, ZN => VGA_l072_n_233);
  VGA_l072_g12414 : OAI211D0BWP7T port map(A1 => VGA_l072_n_191, A2 => VGA_l072_n_209, B => VGA_l072_n_204, C => VGA_l072_n_199, ZN => VGA_enable6);
  VGA_l072_g12415 : OAI22D0BWP7T port map(A1 => VGA_l072_n_217, A2 => VGA_l072_n_139, B1 => VGA_l072_n_207, B2 => VGA_l072_n_131, ZN => VGA_l072_n_231);
  VGA_l072_g12416 : AOI31D0BWP7T port map(A1 => VGA_l072_n_190, A2 => VGA_l072_n_182, A3 => VGA_l072_n_77, B => VGA_l072_n_229, ZN => VGA_l072_n_230);
  VGA_l072_g12417 : AOI21D0BWP7T port map(A1 => VGA_l072_n_103, A2 => VGA_l072_n_86, B => VGA_l072_n_216, ZN => VGA_l072_n_229);
  VGA_l072_g12418 : AOI31D0BWP7T port map(A1 => VGA_l072_n_145, A2 => VGA_l072_n_88, A3 => VGA_l072_n_75, B => VGA_l072_n_217, ZN => VGA_l072_n_228);
  VGA_l072_g12419 : AOI31D0BWP7T port map(A1 => VGA_l072_n_122, A2 => VGA_l072_n_118, A3 => VGA_l072_n_60, B => VGA_l072_n_214, ZN => VGA_l072_n_227);
  VGA_l072_g12420 : AOI31D0BWP7T port map(A1 => VGA_l072_n_142, A2 => VGA_l072_n_122, A3 => VGA_l072_n_88, B => VGA_l072_n_215, ZN => VGA_l072_n_226);
  VGA_l072_g12421 : AOI22D0BWP7T port map(A1 => VGA_l072_n_205, A2 => VGA_l072_n_195, B1 => VGA_l072_n_119, B2 => VGA_l072_n_89, ZN => VGA_l072_n_225);
  VGA_l072_g12422 : AO21D0BWP7T port map(A1 => VGA_l072_n_123, A2 => VGA_l072_n_91, B => VGA_l072_n_215, Z => VGA_l072_n_224);
  VGA_l072_g12423 : OA21D0BWP7T port map(A1 => VGA_l072_n_208, A2 => VGA_l072_n_157, B => VGA_l072_n_222, Z => VGA_l072_n_223);
  VGA_l072_g12424 : AO31D0BWP7T port map(A1 => VGA_l072_n_135, A2 => VGA_l072_n_68, A3 => VGA_l072_n_69, B => VGA_l072_n_204, Z => VGA_l072_n_222);
  VGA_l072_g12425 : AOI21D0BWP7T port map(A1 => VGA_l072_n_89, A2 => VGA_l072_n_52, B => VGA_l072_n_212, ZN => VGA_l072_n_221);
  VGA_l072_g12426 : AOI31D0BWP7T port map(A1 => VGA_l072_n_132, A2 => VGA_l072_n_76, A3 => VGA_l072_n_58, B => VGA_l072_n_207, ZN => VGA_l072_n_220);
  VGA_l072_g12427 : OA21D0BWP7T port map(A1 => VGA_l072_n_134, A2 => VGA_l072_n_90, B => VGA_l072_n_211, Z => VGA_l072_n_219);
  VGA_l072_g12428 : AOI21D0BWP7T port map(A1 => VGA_l072_n_88, A2 => VGA_l072_n_0, B => VGA_l072_n_204, ZN => VGA_l072_n_218);
  VGA_l072_g12429 : AOI32D0BWP7T port map(A1 => VGA_l072_n_190, A2 => VGA_l072_n_181, A3 => VGA_l072_n_38, B1 => VGA_l072_n_202, B2 => VGA_l072_n_154, ZN => VGA_l072_n_214);
  VGA_l072_g12430 : AOI21D0BWP7T port map(A1 => VGA_l072_n_103, A2 => VGA_l072_n_68, B => VGA_l072_n_208, ZN => VGA_l072_n_213);
  VGA_l072_g12431 : AOI22D0BWP7T port map(A1 => VGA_l072_n_203, A2 => VGA_l072_n_156, B1 => VGA_l072_n_202, B2 => VGA_l072_n_143, ZN => VGA_l072_n_217);
  VGA_l072_g12432 : AOI22D0BWP7T port map(A1 => VGA_l072_n_202, A2 => VGA_l072_n_160, B1 => VGA_l072_n_203, B2 => VGA_l072_n_144, ZN => VGA_l072_n_216);
  VGA_l072_g12433 : AOI32D0BWP7T port map(A1 => VGA_l072_n_198, A2 => VGA_l072_n_1, A3 => VGA_l072_n_104, B1 => VGA_l072_n_203, B2 => VGA_l072_n_155, ZN => VGA_l072_n_215);
  VGA_l072_g12434 : OAI31D0BWP7T port map(A1 => VGA_l072_n_2, A2 => VGA_l072_n_127, A3 => VGA_l072_n_179, B => VGA_l072_n_201, ZN => VGA_l072_n_210);
  VGA_l072_g12435 : NR4D0BWP7T port map(A1 => VGA_l072_n_200, A2 => VGA_l072_n_186, A3 => VGA_l072_n_182, A4 => VGA_l072_n_185, ZN => VGA_l072_n_209);
  VGA_l072_g12436 : MAOI22D0BWP7T port map(A1 => VGA_l072_n_196, A2 => VGA_l072_n_170, B1 => VGA_l072_n_191, B2 => VGA_l072_n_165, ZN => VGA_l072_n_212);
  VGA_l072_g12437 : OAI22D0BWP7T port map(A1 => VGA_l072_n_197, A2 => VGA_l072_n_171, B1 => VGA_l072_n_193, B2 => VGA_l072_n_150, ZN => VGA_l072_n_211);
  VGA_l072_g12438 : CKND1BWP7T port map(I => VGA_l072_n_206, ZN => VGA_l072_n_205);
  VGA_l072_g12439 : AOI22D0BWP7T port map(A1 => VGA_l072_n_196, A2 => VGA_l072_n_169, B1 => VGA_l072_n_194, B2 => VGA_l072_n_151, ZN => VGA_l072_n_208);
  VGA_l072_g12440 : MAOI22D0BWP7T port map(A1 => VGA_l072_n_196, A2 => VGA_l072_n_151, B1 => VGA_l072_n_193, B2 => VGA_l072_n_168, ZN => VGA_l072_n_207);
  VGA_l072_g12441 : OAI22D0BWP7T port map(A1 => VGA_l072_n_197, A2 => VGA_l072_n_167, B1 => VGA_l072_n_191, B2 => VGA_l072_n_176, ZN => VGA_l072_n_206);
  VGA_l072_g12442 : MAOI22D0BWP7T port map(A1 => VGA_l072_n_196, A2 => VGA_l072_n_140, B1 => VGA_l072_n_193, B2 => VGA_l072_n_167, ZN => VGA_l072_n_204);
  VGA_l072_g12443 : INR2D0BWP7T port map(A1 => VGA_l072_n_198, B1 => VGA_l072_n_114, ZN => VGA_l072_n_203);
  VGA_l072_g12444 : INR2D0BWP7T port map(A1 => VGA_l072_n_198, B1 => VGA_l072_n_113, ZN => VGA_l072_n_202);
  VGA_l072_g12445 : CKND1BWP7T port map(I => VGA_l072_n_200, ZN => VGA_l072_n_201);
  VGA_l072_g12446 : OAI21D0BWP7T port map(A1 => VGA_l072_n_177, A2 => VGA_l072_n_161, B => VGA_l072_n_194, ZN => VGA_l072_n_199);
  VGA_l072_g12447 : ND3D0BWP7T port map(A1 => VGA_l072_n_188, A2 => VGA_l072_n_176, A3 => VGA_l072_n_165, ZN => VGA_l072_n_200);
  VGA_l072_g12448 : INVD0BWP7T port map(I => VGA_l072_n_197, ZN => VGA_l072_n_196);
  VGA_l072_g12449 : INR2D0BWP7T port map(A1 => VGA_l072_n_185, B1 => VGA_l072_n_191, ZN => VGA_l072_n_198);
  VGA_l072_g12450 : ND2D0BWP7T port map(A1 => VGA_l072_n_190, A2 => VGA_l072_n_184, ZN => VGA_l072_n_197);
  VGA_l072_g12451 : CKND1BWP7T port map(I => VGA_l072_n_193, ZN => VGA_l072_n_194);
  VGA_l072_g12452 : AOI211D0BWP7T port map(A1 => VGA_l072_n_122, A2 => VGA_l072_n_74, B => VGA_l072_n_191, C => VGA_l072_n_183, ZN => VGA_l072_n_192);
  VGA_l072_g12453 : IND2D0BWP7T port map(A1 => VGA_l072_n_189, B1 => VGA_l072_n_190, ZN => VGA_l072_n_195);
  VGA_l072_g12454 : ND2D0BWP7T port map(A1 => VGA_l072_n_190, A2 => VGA_l072_n_164, ZN => VGA_l072_n_193);
  VGA_l072_g12455 : INVD1BWP7T port map(I => VGA_l072_n_191, ZN => VGA_l072_n_190);
  VGA_l072_g12456 : OAI221D0BWP7T port map(A1 => VGA_l072_n_49, A2 => VGA_l072_n_32, B1 => VGA_l072_n_20, B2 => VGA_l072_n_21, C => VGA_l072_n_187, ZN => VGA_l072_n_191);
  VGA_l072_g12457 : AOI22D0BWP7T port map(A1 => VGA_l072_n_184, A2 => VGA_l072_n_161, B1 => VGA_l072_n_170, B2 => VGA_l072_n_164, ZN => VGA_l072_n_188);
  VGA_l072_g12458 : AOI33D0BWP7T port map(A1 => VGA_l072_n_184, A2 => VGA_l072_n_143, A3 => VGA_l072_n_113, B1 => VGA_l072_n_164, B2 => VGA_l072_n_156, B3 => VGA_l072_n_114, ZN => VGA_l072_n_189);
  VGA_l072_g12459 : AOI211D0BWP7T port map(A1 => VGA_l072_n_173, A2 => VGA_l072_n_136, B => VGA_l072_n_178, C => VGA_l072_n_120, ZN => VGA_l072_n_187);
  VGA_l072_g12460 : OA21D0BWP7T port map(A1 => VGA_l072_n_180, A2 => VGA_l072_n_170, B => VGA_l072_n_184, Z => VGA_l072_n_186);
  VGA_l072_g12461 : NR2D0BWP7T port map(A1 => VGA_l072_n_179, A2 => VGA_l072_n_115, ZN => VGA_l072_n_185);
  VGA_l072_g12462 : NR2D0BWP7T port map(A1 => VGA_l072_n_179, A2 => VGA_l072_n_116, ZN => VGA_l072_n_184);
  VGA_l072_g12463 : CKND1BWP7T port map(I => VGA_l072_n_182, ZN => VGA_l072_n_183);
  VGA_l072_g12464 : AO32D0BWP7T port map(A1 => VGA_l072_n_166, A2 => VGA_l072_n_102, A3 => VGA_l072_n_37, B1 => VGA_l072_n_175, B2 => VGA_y(4), Z => VGA_l072_n_181);
  VGA_l072_g12465 : OAI22D0BWP7T port map(A1 => VGA_l072_n_172, A2 => VGA_l072_n_113, B1 => VGA_l072_n_174, B2 => VGA_l072_n_38, ZN => VGA_l072_n_182);
  VGA_l072_g12466 : IND2D0BWP7T port map(A1 => VGA_l072_n_177, B1 => VGA_l072_n_167, ZN => VGA_l072_n_180);
  VGA_l072_g12467 : MOAI22D0BWP7T port map(A1 => VGA_l072_n_163, A2 => VGA_l072_n_136, B1 => VGA_l072_n_21, B2 => VGA_l072_n_20, ZN => VGA_l072_n_178);
  VGA_l072_g12468 : AOI22D0BWP7T port map(A1 => VGA_l072_n_166, A2 => y_pos_e2(4), B1 => VGA_l072_n_159, B2 => VGA_l072_n_11, ZN => VGA_l072_n_179);
  VGA_l072_g12469 : ND2D0BWP7T port map(A1 => VGA_l072_n_168, A2 => VGA_l072_n_171, ZN => VGA_l072_n_177);
  VGA_l072_g12470 : ND2D0BWP7T port map(A1 => VGA_l072_n_164, A2 => VGA_l072_n_140, ZN => VGA_l072_n_176);
  VGA_l072_g12471 : CKND1BWP7T port map(I => VGA_l072_n_174, ZN => VGA_l072_n_175);
  VGA_l072_g12472 : OAI211D0BWP7T port map(A1 => VGA_l072_n_96, A2 => VGA_l072_n_129, B => VGA_l072_n_153, C => VGA_l072_n_105, ZN => VGA_l072_n_173);
  VGA_l072_g12473 : ND3D0BWP7T port map(A1 => VGA_l072_n_154, A2 => VGA_l072_n_158, A3 => VGA_l072_n_115, ZN => VGA_l072_n_172);
  VGA_l072_g12474 : ND3D0BWP7T port map(A1 => VGA_l072_n_159, A2 => VGA_l072_n_102, A3 => VGA_l072_n_37, ZN => VGA_l072_n_174);
  VGA_l072_g12475 : CKND1BWP7T port map(I => VGA_l072_n_168, ZN => VGA_l072_n_169);
  VGA_l072_g12476 : ND2D0BWP7T port map(A1 => VGA_l072_n_156, A2 => VGA_l072_n_114, ZN => VGA_l072_n_171);
  VGA_l072_g12477 : AN2D1BWP7T port map(A1 => VGA_l072_n_154, A2 => VGA_l072_n_113, Z => VGA_l072_n_170);
  VGA_l072_g12478 : ND2D0BWP7T port map(A1 => VGA_l072_n_160, A2 => VGA_l072_n_113, ZN => VGA_l072_n_168);
  VGA_l072_g12479 : ND2D0BWP7T port map(A1 => VGA_l072_n_155, A2 => VGA_l072_n_114, ZN => VGA_l072_n_167);
  VGA_l072_g12480 : AOI221D0BWP7T port map(A1 => VGA_l072_n_125, A2 => VGA_l072_n_95, B1 => VGA_l072_n_45, B2 => VGA_l072_n_81, C => VGA_l072_n_152, ZN => VGA_l072_n_163);
  VGA_l072_g12481 : AN4D1BWP7T port map(A1 => VGA_l072_n_141, A2 => VGA_l072_n_103, A3 => VGA_l072_n_89, A4 => VGA_l072_n_0, Z => VGA_l072_n_162);
  VGA_l072_g12482 : NR3D0BWP7T port map(A1 => VGA_l072_n_149, A2 => VGA_l072_n_44, A3 => VGA_y(4), ZN => VGA_l072_n_166);
  VGA_l072_g12483 : IND3D0BWP7T port map(A1 => VGA_l072_n_127, B1 => VGA_l072_n_2, B2 => VGA_l072_n_158, ZN => VGA_l072_n_165);
  VGA_l072_g12484 : AN2D1BWP7T port map(A1 => VGA_l072_n_158, A2 => VGA_l072_n_116, Z => VGA_l072_n_164);
  VGA_l072_g12485 : IINR4D0BWP7T port map(A1 => VGA_l072_n_122, A2 => VGA_l072_n_69, B1 => VGA_l072_n_133, B2 => VGA_l072_n_77, ZN => VGA_l072_n_157);
  VGA_l072_g12486 : IND2D0BWP7T port map(A1 => VGA_l072_n_151, B1 => VGA_l072_n_150, ZN => VGA_l072_n_161);
  VGA_l072_g12487 : NR3D0BWP7T port map(A1 => VGA_l072_n_148, A2 => VGA_l072_n_87, A3 => VGA_l072_n_40, ZN => VGA_l072_n_160);
  VGA_l072_g12488 : INR2D0BWP7T port map(A1 => VGA_l072_n_44, B1 => VGA_l072_n_149, ZN => VGA_l072_n_159);
  VGA_l072_g12489 : AOI211D0BWP7T port map(A1 => VGA_l072_n_44, A2 => VGA_l072_n_34, B => VGA_l072_n_149, C => VGA_l072_n_98, ZN => VGA_l072_n_158);
  VGA_l072_g12490 : AOI22D0BWP7T port map(A1 => VGA_l072_n_146, A2 => VGA_l072_n_126, B1 => VGA_l072_n_45, B2 => VGA_l072_n_26, ZN => VGA_l072_n_153);
  VGA_l072_g12491 : OAI22D0BWP7T port map(A1 => VGA_l072_n_146, A2 => VGA_l072_n_130, B1 => VGA_l072_n_97, B2 => VGA_x(5), ZN => VGA_l072_n_152);
  VGA_l072_g12492 : INR3D0BWP7T port map(A1 => VGA_l072_n_148, B1 => VGA_l072_n_40, B2 => VGA_l072_n_87, ZN => VGA_l072_n_156);
  VGA_l072_g12493 : AN3D0BWP7T port map(A1 => VGA_l072_n_147, A2 => VGA_l072_n_87, A3 => VGA_l072_n_39, Z => VGA_l072_n_155);
  VGA_l072_g12494 : INR3D0BWP7T port map(A1 => VGA_l072_n_87, B1 => VGA_l072_n_40, B2 => VGA_l072_n_147, ZN => VGA_l072_n_154);
  VGA_l072_g12495 : AN2D1BWP7T port map(A1 => VGA_l072_n_144, A2 => VGA_l072_n_114, Z => VGA_l072_n_151);
  VGA_l072_g12496 : ND2D0BWP7T port map(A1 => VGA_l072_n_143, A2 => VGA_l072_n_113, ZN => VGA_l072_n_150);
  VGA_l072_g12497 : IND4D0BWP7T port map(A1 => VGA_l072_n_108, B1 => VGA_l072_n_109, B2 => VGA_l072_n_106, B3 => VGA_l072_n_107, ZN => VGA_l072_n_149);
  VGA_l072_g12498 : AN3D0BWP7T port map(A1 => VGA_l072_n_128, A2 => VGA_l072_n_70, A3 => VGA_l072_n_76, Z => VGA_l072_n_145);
  VGA_l072_g12499 : OAI221D0BWP7T port map(A1 => VGA_l072_n_101, A2 => y_pos_e2(1), B1 => VGA_l072_n_4, B2 => VGA_l072_n_82, C => VGA_l072_n_100, ZN => VGA_l072_n_148);
  VGA_l072_g12500 : OAI211D0BWP7T port map(A1 => y_pos_e2(1), A2 => VGA_l072_n_41, B => VGA_l072_n_121, C => VGA_l072_n_101, ZN => VGA_l072_n_147);
  VGA_l072_g12501 : MAOI222D0BWP7T port map(A => VGA_x(2), B => x_pos_e2(2), C => VGA_l072_n_83, ZN => VGA_l072_n_146);
  VGA_l072_g12502 : AN3D0BWP7T port map(A1 => VGA_l072_n_124, A2 => VGA_l072_n_94, A3 => VGA_l072_n_92, Z => VGA_l072_n_142);
  VGA_l072_g12503 : INR3D0BWP7T port map(A1 => VGA_l072_n_128, B1 => VGA_l072_n_72, B2 => VGA_l072_n_77, ZN => VGA_l072_n_141);
  VGA_l072_g12504 : AOI211D0BWP7T port map(A1 => VGA_l072_n_101, A2 => VGA_l072_n_100, B => VGA_l072_n_39, C => VGA_l072_n_43, ZN => VGA_l072_n_144);
  VGA_l072_g12505 : AN4D1BWP7T port map(A1 => VGA_l072_n_101, A2 => VGA_l072_n_100, A3 => VGA_l072_n_42, A4 => VGA_l072_n_40, Z => VGA_l072_n_143);
  VGA_l072_g12506 : INR2D0BWP7T port map(A1 => VGA_l072_n_122, B1 => VGA_l072_n_72, ZN => VGA_l072_n_139);
  VGA_l072_g12507 : AN2D1BWP7T port map(A1 => VGA_l072_n_112, A2 => VGA_l072_n_52, Z => VGA_l072_n_138);
  VGA_l072_g12508 : ND2D0BWP7T port map(A1 => VGA_l072_n_123, A2 => VGA_l072_n_131, ZN => VGA_l072_n_137);
  VGA_l072_g12509 : INR2D0BWP7T port map(A1 => VGA_l072_n_104, B1 => VGA_l072_n_1, ZN => VGA_l072_n_140);
  VGA_l072_g12510 : OA221D0BWP7T port map(A1 => VGA_l072_n_67, A2 => VGA_draw_count6(1), B1 => VGA_l072_n_24, B2 => VGA_l072_n_54, C => VGA_l072_n_74, Z => VGA_l072_n_135);
  VGA_l072_g12511 : OAI211D0BWP7T port map(A1 => VGA_draw_count6(1), A2 => VGA_l072_n_58, B => VGA_l072_n_84, C => VGA_l072_n_74, ZN => VGA_l072_n_134);
  VGA_l072_g12512 : OAI211D0BWP7T port map(A1 => VGA_l072_n_13, A2 => VGA_l072_n_54, B => VGA_l072_n_85, C => VGA_l072_n_75, ZN => VGA_l072_n_133);
  VGA_l072_g12513 : OA21D0BWP7T port map(A1 => VGA_l072_n_14, A2 => VGA_l072_n_3, B => VGA_l072_n_124, Z => VGA_l072_n_132);
  VGA_l072_g12514 : ND2D0BWP7T port map(A1 => VGA_l072_n_110, A2 => VGA_l072_n_105, ZN => VGA_l072_n_136);
  VGA_l072_g12515 : CKND1BWP7T port map(I => VGA_l072_n_129, ZN => VGA_l072_n_130);
  VGA_l072_g12516 : CKND1BWP7T port map(I => VGA_l072_n_125, ZN => VGA_l072_n_126);
  VGA_l072_g12517 : IND2D0BWP7T port map(A1 => VGA_l072_n_100, B1 => y_pos_e2(1), ZN => VGA_l072_n_121);
  VGA_l072_g12518 : MOAI22D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l072_n_10, B1 => VGA_l072_n_49, B2 => VGA_l072_n_32, ZN => VGA_l072_n_120);
  VGA_l072_g12519 : AOI21D0BWP7T port map(A1 => VGA_l072_n_59, A2 => VGA_l072_n_27, B => VGA_l072_n_93, ZN => VGA_l072_n_119);
  VGA_l072_g12520 : AOI211D0BWP7T port map(A1 => VGA_l072_n_55, A2 => VGA_l072_n_24, B => VGA_l072_n_93, C => VGA_l072_n_78, ZN => VGA_l072_n_118);
  VGA_l072_g12521 : OAI221D0BWP7T port map(A1 => VGA_l072_n_62, A2 => VGA_l072_n_0, B1 => VGA_l072_n_29, B2 => VGA_l072_n_64, C => VGA_l072_n_92, ZN => VGA_l072_n_117);
  VGA_l072_g12522 : OA21D0BWP7T port map(A1 => VGA_l072_n_62, A2 => VGA_l072_n_64, B => VGA_l072_n_92, Z => VGA_l072_n_131);
  VGA_l072_g12523 : AOI22D0BWP7T port map(A1 => VGA_l072_n_66, A2 => VGA_l072_n_31, B1 => VGA_l072_n_47, B2 => VGA_x(2), ZN => VGA_l072_n_129);
  VGA_l072_g12524 : NR3D0BWP7T port map(A1 => VGA_l072_n_80, A2 => VGA_l072_n_73, A3 => VGA_l072_n_61, ZN => VGA_l072_n_128);
  VGA_l072_g12525 : IND2D0BWP7T port map(A1 => VGA_l072_n_37, B1 => VGA_l072_n_102, ZN => VGA_l072_n_127);
  VGA_l072_g12526 : OAI22D0BWP7T port map(A1 => VGA_l072_n_66, A2 => VGA_l072_n_31, B1 => VGA_l072_n_47, B2 => VGA_x(2), ZN => VGA_l072_n_125);
  VGA_l072_g12527 : AN3D0BWP7T port map(A1 => VGA_l072_n_68, A2 => VGA_l072_n_75, A3 => VGA_l072_n_69, Z => VGA_l072_n_124);
  VGA_l072_g12528 : AN2D1BWP7T port map(A1 => VGA_l072_n_88, A2 => VGA_l072_n_68, Z => VGA_l072_n_123);
  VGA_l072_g12529 : AN2D1BWP7T port map(A1 => VGA_l072_n_89, A2 => VGA_l072_n_58, Z => VGA_l072_n_122);
  VGA_l072_g12530 : AOI221D0BWP7T port map(A1 => VGA_l072_n_61, A2 => VGA_draw_count6(0), B1 => VGA_l072_n_56, B2 => VGA_l072_n_25, C => VGA_l072_n_80, ZN => VGA_l072_n_112);
  VGA_l072_g12531 : AO222D0BWP7T port map(A1 => VGA_l072_n_61, A2 => VGA_l072_n_24, B1 => VGA_l072_n_55, B2 => VGA_l072_n_13, C1 => VGA_l072_n_53, C2 => VGA_l072_n_27, Z => VGA_l072_n_111);
  VGA_l072_g12532 : OAI22D0BWP7T port map(A1 => VGA_l072_n_45, A2 => VGA_l072_n_26, B1 => VGA_l072_n_46, B2 => VGA_l072_n_16, ZN => VGA_l072_n_110);
  VGA_l072_g12533 : MAOI22D0BWP7T port map(A1 => VGA_l072_n_50, A2 => VGA_l072_n_35, B1 => VGA_l072_n_50, B2 => VGA_l072_n_35, ZN => VGA_l072_n_109);
  VGA_l072_g12534 : OAI22D0BWP7T port map(A1 => VGA_l072_n_65, A2 => VGA_l072_n_15, B1 => VGA_l072_n_36, B2 => VGA_y(9), ZN => VGA_l072_n_108);
  VGA_l072_g12535 : AOI22D0BWP7T port map(A1 => VGA_l072_n_65, A2 => VGA_l072_n_15, B1 => VGA_l072_n_36, B2 => VGA_y(9), ZN => VGA_l072_n_107);
  VGA_l072_g12536 : MAOI22D0BWP7T port map(A1 => VGA_l072_n_48, A2 => VGA_l072_n_28, B1 => VGA_l072_n_48, B2 => VGA_l072_n_28, ZN => VGA_l072_n_106);
  VGA_l072_g12538 : MAOI22D0BWP7T port map(A1 => VGA_l072_n_38, A2 => VGA_l072_n_19, B1 => VGA_l072_n_38, B2 => VGA_l072_n_19, ZN => VGA_l072_n_116);
  VGA_l072_g12540 : MOAI22D0BWP7T port map(A1 => VGA_l072_n_38, A2 => VGA_l072_n_22, B1 => VGA_l072_n_38, B2 => VGA_l072_n_22, ZN => VGA_l072_n_115);
  VGA_l072_g12541 : MAOI22D0BWP7T port map(A1 => VGA_l072_n_37, A2 => VGA_l072_n_33, B1 => VGA_l072_n_37, B2 => VGA_l072_n_33, ZN => VGA_l072_n_114);
  VGA_l072_g12542 : MOAI22D0BWP7T port map(A1 => VGA_l072_n_37, A2 => VGA_l072_n_23, B1 => VGA_l072_n_37, B2 => VGA_l072_n_23, ZN => VGA_l072_n_113);
  VGA_l072_g12543 : AOI21D0BWP7T port map(A1 => VGA_l072_n_56, A2 => VGA_l072_n_24, B => VGA_l072_n_63, ZN => VGA_l072_n_99);
  VGA_l072_g12544 : NR2D0BWP7T port map(A1 => VGA_l072_n_44, A2 => VGA_l072_n_34, ZN => VGA_l072_n_98);
  VGA_l072_g12545 : IND2D0BWP7T port map(A1 => VGA_l072_n_46, B1 => x_pos_e2(5), ZN => VGA_l072_n_97);
  VGA_l072_g12546 : ND2D0BWP7T port map(A1 => VGA_l072_n_46, A2 => VGA_l072_n_16, ZN => VGA_l072_n_105);
  VGA_l072_g12547 : NR2D0BWP7T port map(A1 => VGA_l072_n_66, A2 => VGA_l072_n_31, ZN => VGA_l072_n_96);
  VGA_l072_g12548 : NR2D0BWP7T port map(A1 => VGA_l072_n_71, A2 => VGA_l072_n_41, ZN => VGA_l072_n_104);
  VGA_l072_g12550 : NR2D0BWP7T port map(A1 => VGA_l072_n_79, A2 => VGA_l072_n_78, ZN => VGA_l072_n_103);
  VGA_l072_g12551 : NR2D0BWP7T port map(A1 => VGA_l072_n_71, A2 => VGA_l072_n_82, ZN => VGA_l072_n_102);
  VGA_l072_g12552 : ND2D0BWP7T port map(A1 => VGA_l072_n_82, A2 => VGA_y(1), ZN => VGA_l072_n_101);
  VGA_l072_g12553 : IND2D0BWP7T port map(A1 => VGA_y(1), B1 => VGA_l072_n_41, ZN => VGA_l072_n_100);
  VGA_l072_g12554 : CKND1BWP7T port map(I => VGA_l072_n_90, ZN => VGA_l072_n_91);
  VGA_l072_g12555 : AOI21D0BWP7T port map(A1 => VGA_l072_n_59, A2 => VGA_l072_n_25, B => VGA_l072_n_73, ZN => VGA_l072_n_86);
  VGA_l072_g12556 : OAI21D0BWP7T port map(A1 => VGA_l072_n_56, A2 => VGA_l072_n_53, B => VGA_l072_n_24, ZN => VGA_l072_n_85);
  VGA_l072_g12557 : AO21D0BWP7T port map(A1 => VGA_l072_n_60, A2 => VGA_l072_n_54, B => VGA_l072_n_62, Z => VGA_l072_n_84);
  VGA_l072_g12558 : IAO21D0BWP7T port map(A1 => VGA_l072_n_60, A2 => VGA_l072_n_13, B => VGA_l072_n_55, ZN => VGA_l072_n_94);
  VGA_l072_g12559 : OAI21D0BWP7T port map(A1 => VGA_l072_n_52, A2 => VGA_draw_count6(1), B => VGA_l072_n_70, ZN => VGA_l072_n_93);
  VGA_l072_g12560 : AOI22D0BWP7T port map(A1 => VGA_l072_n_51, A2 => VGA_x(0), B1 => VGA_x(1), B2 => VGA_l072_n_6, ZN => VGA_l072_n_83);
  VGA_l072_g12561 : OA22D0BWP7T port map(A1 => VGA_l072_n_64, A2 => VGA_l072_n_12, B1 => VGA_l072_n_25, B2 => VGA_l072_n_0, Z => VGA_l072_n_92);
  VGA_l072_g12562 : OAI21D0BWP7T port map(A1 => VGA_l072_n_57, A2 => VGA_l072_n_13, B => VGA_l072_n_69, ZN => VGA_l072_n_90);
  VGA_l072_g12563 : AOI22D0BWP7T port map(A1 => VGA_l072_n_56, A2 => VGA_l072_n_13, B1 => VGA_l072_n_59, B2 => VGA_l072_n_24, ZN => VGA_l072_n_89);
  VGA_l072_g12564 : IAO21D0BWP7T port map(A1 => VGA_l072_n_0, A2 => VGA_l072_n_24, B => VGA_l072_n_79, ZN => VGA_l072_n_88);
  VGA_l072_g12565 : MOAI22D0BWP7T port map(A1 => VGA_l072_n_43, A2 => VGA_y(0), B1 => VGA_l072_n_43, B2 => VGA_y(0), ZN => VGA_l072_n_87);
  VGA_l072_g12568 : INVD0BWP7T port map(I => VGA_l072_n_41, ZN => VGA_l072_n_82);
  VGA_l072_g12569 : CKND1BWP7T port map(I => VGA_l072_n_26, ZN => VGA_l072_n_81);
  VGA_l072_g12570 : NR2D0BWP7T port map(A1 => VGA_l072_n_54, A2 => VGA_draw_count6(1), ZN => VGA_l072_n_80);
  VGA_l072_g12571 : INR2D0BWP7T port map(A1 => VGA_l072_n_63, B1 => VGA_l072_n_25, ZN => VGA_l072_n_79);
  VGA_l072_g12572 : NR2D0BWP7T port map(A1 => VGA_l072_n_0, A2 => VGA_draw_count6(1), ZN => VGA_l072_n_78);
  VGA_l072_g12573 : NR2D0BWP7T port map(A1 => VGA_l072_n_57, A2 => VGA_l072_n_29, ZN => VGA_l072_n_77);
  VGA_l072_g12574 : ND2D0BWP7T port map(A1 => VGA_l072_n_55, A2 => VGA_draw_count6(1), ZN => VGA_l072_n_76);
  VGA_l072_g12575 : ND2D0BWP7T port map(A1 => VGA_l072_n_53, A2 => VGA_l072_n_13, ZN => VGA_l072_n_75);
  VGA_l072_g12576 : ND2D0BWP7T port map(A1 => VGA_l072_n_53, A2 => VGA_draw_count6(1), ZN => VGA_l072_n_74);
  VGA_l072_g12577 : NR2D0BWP7T port map(A1 => VGA_l072_n_56, A2 => VGA_l072_n_59, ZN => VGA_l072_n_67);
  VGA_l072_g12578 : AN2D1BWP7T port map(A1 => VGA_l072_n_63, A2 => VGA_l072_n_27, Z => VGA_l072_n_73);
  VGA_l072_g12579 : NR2D0BWP7T port map(A1 => VGA_l072_n_52, A2 => VGA_l072_n_13, ZN => VGA_l072_n_72);
  VGA_l072_g12580 : ND2D0BWP7T port map(A1 => VGA_l072_n_40, A2 => VGA_l072_n_43, ZN => VGA_l072_n_71);
  VGA_l072_g12581 : IND2D0BWP7T port map(A1 => VGA_l072_n_62, B1 => VGA_l072_n_56, ZN => VGA_l072_n_70);
  VGA_l072_g12582 : ND2D0BWP7T port map(A1 => VGA_l072_n_63, A2 => VGA_l072_n_13, ZN => VGA_l072_n_69);
  VGA_l072_g12583 : IND2D0BWP7T port map(A1 => VGA_l072_n_62, B1 => VGA_l072_n_63, ZN => VGA_l072_n_68);
  VGA_l072_g12584 : INVD0BWP7T port map(I => VGA_l072_n_61, ZN => VGA_l072_n_60);
  VGA_l072_g12585 : INVD0BWP7T port map(I => VGA_l072_n_59, ZN => VGA_l072_n_58);
  VGA_l072_g12586 : INVD1BWP7T port map(I => VGA_l072_n_57, ZN => VGA_l072_n_56);
  VGA_l072_g12587 : INVD0BWP7T port map(I => VGA_l072_n_55, ZN => VGA_l072_n_54);
  VGA_l072_g12588 : INVD0BWP7T port map(I => VGA_l072_n_53, ZN => VGA_l072_n_52);
  VGA_l072_g12589 : IAO21D0BWP7T port map(A1 => VGA_x(1), A2 => VGA_l072_n_6, B => x_pos_e2(0), ZN => VGA_l072_n_51);
  VGA_l072_g12590 : OAI21D0BWP7T port map(A1 => VGA_l072_n_7, A2 => x_pos_e2(4), B => VGA_l072_n_26, ZN => VGA_l072_n_66);
  VGA_l072_g12591 : AOI21D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l072_n_5, B => VGA_l072_n_28, ZN => VGA_l072_n_65);
  VGA_l072_g12592 : IND2D0BWP7T port map(A1 => VGA_l072_n_30, B1 => VGA_draw_count6(4), ZN => VGA_l072_n_64);
  VGA_l072_g12593 : INR2D0BWP7T port map(A1 => VGA_draw_count6(4), B1 => VGA_l072_n_17, ZN => VGA_l072_n_63);
  VGA_l072_g12594 : INR2D0BWP7T port map(A1 => VGA_l072_n_29, B1 => VGA_l072_n_27, ZN => VGA_l072_n_62);
  VGA_l072_g12596 : NR2D0BWP7T port map(A1 => VGA_l072_n_14, A2 => VGA_draw_count6(4), ZN => VGA_l072_n_61);
  VGA_l072_g12597 : NR2D0BWP7T port map(A1 => VGA_l072_n_30, A2 => VGA_draw_count6(4), ZN => VGA_l072_n_59);
  VGA_l072_g12598 : IND2D0BWP7T port map(A1 => VGA_l072_n_14, B1 => VGA_draw_count6(4), ZN => VGA_l072_n_57);
  VGA_l072_g12599 : NR2D0BWP7T port map(A1 => VGA_l072_n_17, A2 => VGA_draw_count6(4), ZN => VGA_l072_n_55);
  VGA_l072_g12600 : NR2D0BWP7T port map(A1 => VGA_l072_n_18, A2 => VGA_draw_count6(4), ZN => VGA_l072_n_53);
  VGA_l072_g12601 : CKND1BWP7T port map(I => VGA_l072_n_43, ZN => VGA_l072_n_42);
  VGA_l072_g12602 : CKND1BWP7T port map(I => VGA_l072_n_40, ZN => VGA_l072_n_39);
  VGA_l072_g12603 : MOAI22D0BWP7T port map(A1 => VGA_y(8), A2 => y_pos_e2(8), B1 => VGA_y(8), B2 => y_pos_e2(8), ZN => VGA_l072_n_50);
  VGA_l072_g12604 : MOAI22D0BWP7T port map(A1 => VGA_x(7), A2 => x_pos_e2(7), B1 => VGA_x(7), B2 => x_pos_e2(7), ZN => VGA_l072_n_49);
  VGA_l072_g12605 : MOAI22D0BWP7T port map(A1 => VGA_y(7), A2 => y_pos_e2(7), B1 => VGA_y(7), B2 => y_pos_e2(7), ZN => VGA_l072_n_48);
  VGA_l072_g12606 : MAOI22D0BWP7T port map(A1 => VGA_x(3), A2 => x_pos_e2(3), B1 => VGA_x(3), B2 => x_pos_e2(3), ZN => VGA_l072_n_47);
  VGA_l072_g12607 : MOAI22D0BWP7T port map(A1 => VGA_x(6), A2 => x_pos_e2(6), B1 => VGA_x(6), B2 => x_pos_e2(6), ZN => VGA_l072_n_46);
  VGA_l072_g12608 : MOAI22D0BWP7T port map(A1 => VGA_x(5), A2 => x_pos_e2(5), B1 => VGA_x(5), B2 => x_pos_e2(5), ZN => VGA_l072_n_45);
  VGA_l072_g12609 : MAOI22D0BWP7T port map(A1 => VGA_y(5), A2 => y_pos_e2(5), B1 => VGA_y(5), B2 => y_pos_e2(5), ZN => VGA_l072_n_44);
  VGA_l072_g12610 : MOAI22D0BWP7T port map(A1 => VGA_y(1), A2 => y_pos_e2(1), B1 => VGA_y(1), B2 => y_pos_e2(1), ZN => VGA_l072_n_43);
  VGA_l072_g12611 : MOAI22D0BWP7T port map(A1 => VGA_y(2), A2 => y_pos_e2(2), B1 => VGA_y(2), B2 => y_pos_e2(2), ZN => VGA_l072_n_41);
  VGA_l072_g12612 : MOAI22D0BWP7T port map(A1 => VGA_y(0), A2 => y_pos_e2(0), B1 => VGA_y(0), B2 => y_pos_e2(0), ZN => VGA_l072_n_40);
  VGA_l072_g12613 : MAOI22D0BWP7T port map(A1 => VGA_y(4), A2 => y_pos_e2(4), B1 => VGA_y(4), B2 => y_pos_e2(4), ZN => VGA_l072_n_38);
  VGA_l072_g12614 : MOAI22D0BWP7T port map(A1 => VGA_y(3), A2 => y_pos_e2(3), B1 => VGA_y(3), B2 => y_pos_e2(3), ZN => VGA_l072_n_37);
  VGA_l072_g12615 : INVD1BWP7T port map(I => VGA_l072_n_25, ZN => VGA_l072_n_24);
  VGA_l072_g12616 : IND2D0BWP7T port map(A1 => VGA_y(8), B1 => y_pos_e2(8), ZN => VGA_l072_n_36);
  VGA_l072_g12617 : INR2D0BWP7T port map(A1 => y_pos_e2(7), B1 => VGA_y(7), ZN => VGA_l072_n_35);
  VGA_l072_g12618 : IND2D0BWP7T port map(A1 => y_pos_e2(4), B1 => VGA_y(4), ZN => VGA_l072_n_34);
  VGA_l072_g12619 : IND2D0BWP7T port map(A1 => y_pos_e2(2), B1 => VGA_y(2), ZN => VGA_l072_n_33);
  VGA_l072_g12620 : IND2D0BWP7T port map(A1 => x_pos_e2(6), B1 => VGA_x(6), ZN => VGA_l072_n_32);
  VGA_l072_g12621 : IND2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_e2(3), ZN => VGA_l072_n_31);
  VGA_l072_g12622 : ND2D0BWP7T port map(A1 => VGA_draw_count6(2), A2 => VGA_draw_count6(3), ZN => VGA_l072_n_30);
  VGA_l072_g12623 : ND2D0BWP7T port map(A1 => VGA_l072_n_3, A2 => VGA_draw_count6(0), ZN => VGA_l072_n_29);
  VGA_l072_g12624 : NR2D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l072_n_5, ZN => VGA_l072_n_28);
  VGA_l072_g12625 : NR2D0BWP7T port map(A1 => VGA_l072_n_3, A2 => VGA_draw_count6(0), ZN => VGA_l072_n_27);
  VGA_l072_g12626 : ND2D0BWP7T port map(A1 => VGA_l072_n_7, A2 => x_pos_e2(4), ZN => VGA_l072_n_26);
  VGA_l072_g12627 : ND2D0BWP7T port map(A1 => VGA_draw_count6(1), A2 => VGA_draw_count6(0), ZN => VGA_l072_n_25);
  VGA_l072_g12629 : CKND1BWP7T port map(I => VGA_l072_n_13, ZN => VGA_l072_n_12);
  VGA_l072_g12630 : IND2D0BWP7T port map(A1 => VGA_y(4), B1 => y_pos_e2(4), ZN => VGA_l072_n_11);
  VGA_l072_g12631 : ND2D0BWP7T port map(A1 => VGA_l072_n_8, A2 => y_pos_e2(2), ZN => VGA_l072_n_23);
  VGA_l072_g12632 : NR2D0BWP7T port map(A1 => VGA_l072_n_9, A2 => y_pos_e2(3), ZN => VGA_l072_n_22);
  VGA_l072_g12633 : INR2D0BWP7T port map(A1 => x_pos_e2(7), B1 => VGA_x(7), ZN => VGA_l072_n_21);
  VGA_l072_g12634 : ND2D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l072_n_10, ZN => VGA_l072_n_20);
  VGA_l072_g12635 : INR2D0BWP7T port map(A1 => y_pos_e2(3), B1 => VGA_y(3), ZN => VGA_l072_n_19);
  VGA_l072_g12636 : IND2D0BWP7T port map(A1 => VGA_draw_count6(2), B1 => VGA_draw_count6(3), ZN => VGA_l072_n_18);
  VGA_l072_g12637 : IND2D0BWP7T port map(A1 => VGA_draw_count6(3), B1 => VGA_draw_count6(2), ZN => VGA_l072_n_17);
  VGA_l072_g12638 : INR2D0BWP7T port map(A1 => VGA_x(5), B1 => x_pos_e2(5), ZN => VGA_l072_n_16);
  VGA_l072_g12639 : IND2D0BWP7T port map(A1 => y_pos_e2(5), B1 => VGA_y(5), ZN => VGA_l072_n_15);
  VGA_l072_g12640 : OR2D0BWP7T port map(A1 => VGA_draw_count6(2), A2 => VGA_draw_count6(3), Z => VGA_l072_n_14);
  VGA_l072_g12641 : NR2D0BWP7T port map(A1 => VGA_draw_count6(1), A2 => VGA_draw_count6(0), ZN => VGA_l072_n_13);
  VGA_l072_g12642 : CKND1BWP7T port map(I => x_pos_e2(8), ZN => VGA_l072_n_10);
  VGA_l072_g12643 : CKND1BWP7T port map(I => VGA_y(3), ZN => VGA_l072_n_9);
  VGA_l072_g12644 : CKND1BWP7T port map(I => VGA_y(2), ZN => VGA_l072_n_8);
  VGA_l072_g12645 : CKND1BWP7T port map(I => VGA_x(4), ZN => VGA_l072_n_7);
  VGA_l072_g12646 : CKND1BWP7T port map(I => x_pos_e2(1), ZN => VGA_l072_n_6);
  VGA_l072_g12647 : CKND1BWP7T port map(I => y_pos_e2(6), ZN => VGA_l072_n_5);
  VGA_l072_g12648 : CKND1BWP7T port map(I => y_pos_e2(1), ZN => VGA_l072_n_4);
  VGA_l072_g12649 : INVD0BWP7T port map(I => VGA_draw_count6(1), ZN => VGA_l072_n_3);
  VGA_l072_g2 : MUX2ND0BWP7T port map(I0 => VGA_y(3), I1 => VGA_l072_n_9, S => VGA_l072_n_38, ZN => VGA_l072_n_2);
  VGA_l072_g12650 : MUX2ND0BWP7T port map(I0 => VGA_l072_n_8, I1 => VGA_y(2), S => VGA_l072_n_37, ZN => VGA_l072_n_1);
  VGA_l072_g12651 : IND2D1BWP7T port map(A1 => VGA_l072_n_18, B1 => VGA_draw_count6(4), ZN => VGA_l072_n_0);
  VGA_l072_g12652 : INVD0BWP7T port map(I => VGA_l072_n_66, ZN => VGA_l072_n_95);
  VGA_l073_g12402 : OAI211D0BWP7T port map(A1 => VGA_l073_n_76, A2 => VGA_l073_n_195, B => VGA_l073_n_243, C => VGA_l073_n_223, ZN => VGA_r7);
  VGA_l073_g12403 : AOI211D0BWP7T port map(A1 => VGA_l073_n_206, A2 => VGA_l073_n_111, B => VGA_l073_n_242, C => VGA_l073_n_225, ZN => VGA_l073_n_243);
  VGA_l073_g12404 : OAI211D0BWP7T port map(A1 => VGA_l073_n_162, A2 => VGA_l073_n_216, B => VGA_l073_n_241, C => VGA_l073_n_238, ZN => VGA_l073_n_242);
  VGA_l073_g12405 : NR4D0BWP7T port map(A1 => VGA_l073_n_239, A2 => VGA_l073_n_227, A3 => VGA_l073_n_219, A4 => VGA_l073_n_220, ZN => VGA_l073_n_241);
  VGA_l073_g12406 : OAI211D0BWP7T port map(A1 => VGA_l073_n_91, A2 => VGA_l073_n_212, B => VGA_l073_n_237, C => VGA_l073_n_235, ZN => VGA_g7);
  VGA_l073_g12407 : NR4D0BWP7T port map(A1 => VGA_l073_n_233, A2 => VGA_l073_n_191, A3 => VGA_l073_n_151, A4 => VGA_l073_n_138, ZN => VGA_l073_n_239);
  VGA_l073_g12408 : NR4D0BWP7T port map(A1 => VGA_l073_n_226, A2 => VGA_l073_n_228, A3 => VGA_l073_n_221, A4 => VGA_l073_n_192, ZN => VGA_l073_n_238);
  VGA_l073_g12409 : AOI211D0BWP7T port map(A1 => VGA_l073_n_206, A2 => VGA_l073_n_117, B => VGA_l073_n_236, C => VGA_l073_n_218, ZN => VGA_l073_n_237);
  VGA_l073_g12410 : OAI211D0BWP7T port map(A1 => VGA_l073_n_99, A2 => VGA_l073_n_195, B => VGA_l073_n_230, C => VGA_l073_n_224, ZN => VGA_l073_n_236);
  VGA_l073_g12411 : AOI211D0BWP7T port map(A1 => VGA_l073_n_211, A2 => VGA_l073_n_137, B => VGA_l073_n_231, C => VGA_l073_n_213, ZN => VGA_l073_n_235);
  VGA_l073_g12412 : OAI32D0BWP7T port map(A1 => VGA_l073_n_24, A2 => VGA_l073_n_60, A3 => VGA_l073_n_216, B1 => VGA_l073_n_94, B2 => VGA_l073_n_215, ZN => VGA_b7);
  VGA_l073_g12413 : ND4D0BWP7T port map(A1 => VGA_l073_n_210, A2 => VGA_l073_n_189, A3 => VGA_l073_n_176, A4 => VGA_l073_n_165, ZN => VGA_l073_n_233);
  VGA_l073_g12414 : OAI211D0BWP7T port map(A1 => VGA_l073_n_191, A2 => VGA_l073_n_209, B => VGA_l073_n_204, C => VGA_l073_n_199, ZN => VGA_enable7);
  VGA_l073_g12415 : OAI22D0BWP7T port map(A1 => VGA_l073_n_217, A2 => VGA_l073_n_139, B1 => VGA_l073_n_207, B2 => VGA_l073_n_131, ZN => VGA_l073_n_231);
  VGA_l073_g12416 : AOI31D0BWP7T port map(A1 => VGA_l073_n_190, A2 => VGA_l073_n_182, A3 => VGA_l073_n_77, B => VGA_l073_n_229, ZN => VGA_l073_n_230);
  VGA_l073_g12417 : AOI21D0BWP7T port map(A1 => VGA_l073_n_103, A2 => VGA_l073_n_86, B => VGA_l073_n_216, ZN => VGA_l073_n_229);
  VGA_l073_g12418 : AOI31D0BWP7T port map(A1 => VGA_l073_n_145, A2 => VGA_l073_n_88, A3 => VGA_l073_n_75, B => VGA_l073_n_217, ZN => VGA_l073_n_228);
  VGA_l073_g12419 : AOI31D0BWP7T port map(A1 => VGA_l073_n_122, A2 => VGA_l073_n_118, A3 => VGA_l073_n_60, B => VGA_l073_n_214, ZN => VGA_l073_n_227);
  VGA_l073_g12420 : AOI31D0BWP7T port map(A1 => VGA_l073_n_142, A2 => VGA_l073_n_122, A3 => VGA_l073_n_88, B => VGA_l073_n_215, ZN => VGA_l073_n_226);
  VGA_l073_g12421 : AOI22D0BWP7T port map(A1 => VGA_l073_n_205, A2 => VGA_l073_n_195, B1 => VGA_l073_n_119, B2 => VGA_l073_n_89, ZN => VGA_l073_n_225);
  VGA_l073_g12422 : AO21D0BWP7T port map(A1 => VGA_l073_n_123, A2 => VGA_l073_n_91, B => VGA_l073_n_215, Z => VGA_l073_n_224);
  VGA_l073_g12423 : OA21D0BWP7T port map(A1 => VGA_l073_n_208, A2 => VGA_l073_n_157, B => VGA_l073_n_222, Z => VGA_l073_n_223);
  VGA_l073_g12424 : AO31D0BWP7T port map(A1 => VGA_l073_n_135, A2 => VGA_l073_n_68, A3 => VGA_l073_n_69, B => VGA_l073_n_204, Z => VGA_l073_n_222);
  VGA_l073_g12425 : AOI21D0BWP7T port map(A1 => VGA_l073_n_89, A2 => VGA_l073_n_52, B => VGA_l073_n_212, ZN => VGA_l073_n_221);
  VGA_l073_g12426 : AOI31D0BWP7T port map(A1 => VGA_l073_n_132, A2 => VGA_l073_n_76, A3 => VGA_l073_n_58, B => VGA_l073_n_207, ZN => VGA_l073_n_220);
  VGA_l073_g12427 : OA21D0BWP7T port map(A1 => VGA_l073_n_134, A2 => VGA_l073_n_90, B => VGA_l073_n_211, Z => VGA_l073_n_219);
  VGA_l073_g12428 : AOI21D0BWP7T port map(A1 => VGA_l073_n_88, A2 => VGA_l073_n_0, B => VGA_l073_n_204, ZN => VGA_l073_n_218);
  VGA_l073_g12429 : AOI32D0BWP7T port map(A1 => VGA_l073_n_190, A2 => VGA_l073_n_181, A3 => VGA_l073_n_38, B1 => VGA_l073_n_202, B2 => VGA_l073_n_154, ZN => VGA_l073_n_214);
  VGA_l073_g12430 : AOI21D0BWP7T port map(A1 => VGA_l073_n_103, A2 => VGA_l073_n_68, B => VGA_l073_n_208, ZN => VGA_l073_n_213);
  VGA_l073_g12431 : AOI22D0BWP7T port map(A1 => VGA_l073_n_203, A2 => VGA_l073_n_156, B1 => VGA_l073_n_202, B2 => VGA_l073_n_143, ZN => VGA_l073_n_217);
  VGA_l073_g12432 : AOI22D0BWP7T port map(A1 => VGA_l073_n_202, A2 => VGA_l073_n_160, B1 => VGA_l073_n_203, B2 => VGA_l073_n_144, ZN => VGA_l073_n_216);
  VGA_l073_g12433 : AOI32D0BWP7T port map(A1 => VGA_l073_n_198, A2 => VGA_l073_n_1, A3 => VGA_l073_n_104, B1 => VGA_l073_n_203, B2 => VGA_l073_n_155, ZN => VGA_l073_n_215);
  VGA_l073_g12434 : OAI31D0BWP7T port map(A1 => VGA_l073_n_2, A2 => VGA_l073_n_127, A3 => VGA_l073_n_179, B => VGA_l073_n_201, ZN => VGA_l073_n_210);
  VGA_l073_g12435 : NR4D0BWP7T port map(A1 => VGA_l073_n_200, A2 => VGA_l073_n_186, A3 => VGA_l073_n_182, A4 => VGA_l073_n_185, ZN => VGA_l073_n_209);
  VGA_l073_g12436 : MAOI22D0BWP7T port map(A1 => VGA_l073_n_196, A2 => VGA_l073_n_170, B1 => VGA_l073_n_191, B2 => VGA_l073_n_165, ZN => VGA_l073_n_212);
  VGA_l073_g12437 : OAI22D0BWP7T port map(A1 => VGA_l073_n_197, A2 => VGA_l073_n_171, B1 => VGA_l073_n_193, B2 => VGA_l073_n_150, ZN => VGA_l073_n_211);
  VGA_l073_g12438 : CKND1BWP7T port map(I => VGA_l073_n_206, ZN => VGA_l073_n_205);
  VGA_l073_g12439 : AOI22D0BWP7T port map(A1 => VGA_l073_n_196, A2 => VGA_l073_n_169, B1 => VGA_l073_n_194, B2 => VGA_l073_n_151, ZN => VGA_l073_n_208);
  VGA_l073_g12440 : MAOI22D0BWP7T port map(A1 => VGA_l073_n_196, A2 => VGA_l073_n_151, B1 => VGA_l073_n_193, B2 => VGA_l073_n_168, ZN => VGA_l073_n_207);
  VGA_l073_g12441 : OAI22D0BWP7T port map(A1 => VGA_l073_n_197, A2 => VGA_l073_n_167, B1 => VGA_l073_n_191, B2 => VGA_l073_n_176, ZN => VGA_l073_n_206);
  VGA_l073_g12442 : MAOI22D0BWP7T port map(A1 => VGA_l073_n_196, A2 => VGA_l073_n_140, B1 => VGA_l073_n_193, B2 => VGA_l073_n_167, ZN => VGA_l073_n_204);
  VGA_l073_g12443 : INR2D0BWP7T port map(A1 => VGA_l073_n_198, B1 => VGA_l073_n_114, ZN => VGA_l073_n_203);
  VGA_l073_g12444 : INR2D0BWP7T port map(A1 => VGA_l073_n_198, B1 => VGA_l073_n_113, ZN => VGA_l073_n_202);
  VGA_l073_g12445 : CKND1BWP7T port map(I => VGA_l073_n_200, ZN => VGA_l073_n_201);
  VGA_l073_g12446 : OAI21D0BWP7T port map(A1 => VGA_l073_n_177, A2 => VGA_l073_n_161, B => VGA_l073_n_194, ZN => VGA_l073_n_199);
  VGA_l073_g12447 : ND3D0BWP7T port map(A1 => VGA_l073_n_188, A2 => VGA_l073_n_176, A3 => VGA_l073_n_165, ZN => VGA_l073_n_200);
  VGA_l073_g12448 : INVD0BWP7T port map(I => VGA_l073_n_197, ZN => VGA_l073_n_196);
  VGA_l073_g12449 : INR2D0BWP7T port map(A1 => VGA_l073_n_185, B1 => VGA_l073_n_191, ZN => VGA_l073_n_198);
  VGA_l073_g12450 : ND2D0BWP7T port map(A1 => VGA_l073_n_190, A2 => VGA_l073_n_184, ZN => VGA_l073_n_197);
  VGA_l073_g12451 : CKND1BWP7T port map(I => VGA_l073_n_193, ZN => VGA_l073_n_194);
  VGA_l073_g12452 : AOI211D0BWP7T port map(A1 => VGA_l073_n_122, A2 => VGA_l073_n_74, B => VGA_l073_n_191, C => VGA_l073_n_183, ZN => VGA_l073_n_192);
  VGA_l073_g12453 : IND2D0BWP7T port map(A1 => VGA_l073_n_189, B1 => VGA_l073_n_190, ZN => VGA_l073_n_195);
  VGA_l073_g12454 : ND2D0BWP7T port map(A1 => VGA_l073_n_190, A2 => VGA_l073_n_164, ZN => VGA_l073_n_193);
  VGA_l073_g12455 : INVD1BWP7T port map(I => VGA_l073_n_191, ZN => VGA_l073_n_190);
  VGA_l073_g12456 : OAI221D0BWP7T port map(A1 => VGA_l073_n_49, A2 => VGA_l073_n_32, B1 => VGA_l073_n_20, B2 => VGA_l073_n_21, C => VGA_l073_n_187, ZN => VGA_l073_n_191);
  VGA_l073_g12457 : AOI22D0BWP7T port map(A1 => VGA_l073_n_184, A2 => VGA_l073_n_161, B1 => VGA_l073_n_170, B2 => VGA_l073_n_164, ZN => VGA_l073_n_188);
  VGA_l073_g12458 : AOI33D0BWP7T port map(A1 => VGA_l073_n_184, A2 => VGA_l073_n_143, A3 => VGA_l073_n_113, B1 => VGA_l073_n_164, B2 => VGA_l073_n_156, B3 => VGA_l073_n_114, ZN => VGA_l073_n_189);
  VGA_l073_g12459 : AOI211D0BWP7T port map(A1 => VGA_l073_n_173, A2 => VGA_l073_n_136, B => VGA_l073_n_178, C => VGA_l073_n_120, ZN => VGA_l073_n_187);
  VGA_l073_g12460 : OA21D0BWP7T port map(A1 => VGA_l073_n_180, A2 => VGA_l073_n_170, B => VGA_l073_n_184, Z => VGA_l073_n_186);
  VGA_l073_g12461 : NR2D0BWP7T port map(A1 => VGA_l073_n_179, A2 => VGA_l073_n_115, ZN => VGA_l073_n_185);
  VGA_l073_g12462 : NR2D0BWP7T port map(A1 => VGA_l073_n_179, A2 => VGA_l073_n_116, ZN => VGA_l073_n_184);
  VGA_l073_g12463 : CKND1BWP7T port map(I => VGA_l073_n_182, ZN => VGA_l073_n_183);
  VGA_l073_g12464 : AO32D0BWP7T port map(A1 => VGA_l073_n_166, A2 => VGA_l073_n_102, A3 => VGA_l073_n_37, B1 => VGA_l073_n_175, B2 => VGA_y(4), Z => VGA_l073_n_181);
  VGA_l073_g12465 : OAI22D0BWP7T port map(A1 => VGA_l073_n_172, A2 => VGA_l073_n_113, B1 => VGA_l073_n_174, B2 => VGA_l073_n_38, ZN => VGA_l073_n_182);
  VGA_l073_g12466 : IND2D0BWP7T port map(A1 => VGA_l073_n_177, B1 => VGA_l073_n_167, ZN => VGA_l073_n_180);
  VGA_l073_g12467 : MOAI22D0BWP7T port map(A1 => VGA_l073_n_163, A2 => VGA_l073_n_136, B1 => VGA_l073_n_21, B2 => VGA_l073_n_20, ZN => VGA_l073_n_178);
  VGA_l073_g12468 : AOI22D0BWP7T port map(A1 => VGA_l073_n_166, A2 => y_pos_e3(4), B1 => VGA_l073_n_159, B2 => VGA_l073_n_11, ZN => VGA_l073_n_179);
  VGA_l073_g12469 : ND2D0BWP7T port map(A1 => VGA_l073_n_168, A2 => VGA_l073_n_171, ZN => VGA_l073_n_177);
  VGA_l073_g12470 : ND2D0BWP7T port map(A1 => VGA_l073_n_164, A2 => VGA_l073_n_140, ZN => VGA_l073_n_176);
  VGA_l073_g12471 : CKND1BWP7T port map(I => VGA_l073_n_174, ZN => VGA_l073_n_175);
  VGA_l073_g12472 : OAI211D0BWP7T port map(A1 => VGA_l073_n_96, A2 => VGA_l073_n_129, B => VGA_l073_n_153, C => VGA_l073_n_105, ZN => VGA_l073_n_173);
  VGA_l073_g12473 : ND3D0BWP7T port map(A1 => VGA_l073_n_154, A2 => VGA_l073_n_158, A3 => VGA_l073_n_115, ZN => VGA_l073_n_172);
  VGA_l073_g12474 : ND3D0BWP7T port map(A1 => VGA_l073_n_159, A2 => VGA_l073_n_102, A3 => VGA_l073_n_37, ZN => VGA_l073_n_174);
  VGA_l073_g12475 : CKND1BWP7T port map(I => VGA_l073_n_168, ZN => VGA_l073_n_169);
  VGA_l073_g12476 : ND2D0BWP7T port map(A1 => VGA_l073_n_156, A2 => VGA_l073_n_114, ZN => VGA_l073_n_171);
  VGA_l073_g12477 : AN2D1BWP7T port map(A1 => VGA_l073_n_154, A2 => VGA_l073_n_113, Z => VGA_l073_n_170);
  VGA_l073_g12478 : ND2D0BWP7T port map(A1 => VGA_l073_n_160, A2 => VGA_l073_n_113, ZN => VGA_l073_n_168);
  VGA_l073_g12479 : ND2D0BWP7T port map(A1 => VGA_l073_n_155, A2 => VGA_l073_n_114, ZN => VGA_l073_n_167);
  VGA_l073_g12480 : AOI221D0BWP7T port map(A1 => VGA_l073_n_125, A2 => VGA_l073_n_95, B1 => VGA_l073_n_45, B2 => VGA_l073_n_81, C => VGA_l073_n_152, ZN => VGA_l073_n_163);
  VGA_l073_g12481 : AN4D1BWP7T port map(A1 => VGA_l073_n_141, A2 => VGA_l073_n_103, A3 => VGA_l073_n_89, A4 => VGA_l073_n_0, Z => VGA_l073_n_162);
  VGA_l073_g12482 : NR3D0BWP7T port map(A1 => VGA_l073_n_149, A2 => VGA_l073_n_44, A3 => VGA_y(4), ZN => VGA_l073_n_166);
  VGA_l073_g12483 : IND3D0BWP7T port map(A1 => VGA_l073_n_127, B1 => VGA_l073_n_2, B2 => VGA_l073_n_158, ZN => VGA_l073_n_165);
  VGA_l073_g12484 : AN2D1BWP7T port map(A1 => VGA_l073_n_158, A2 => VGA_l073_n_116, Z => VGA_l073_n_164);
  VGA_l073_g12485 : IINR4D0BWP7T port map(A1 => VGA_l073_n_122, A2 => VGA_l073_n_69, B1 => VGA_l073_n_133, B2 => VGA_l073_n_77, ZN => VGA_l073_n_157);
  VGA_l073_g12486 : IND2D0BWP7T port map(A1 => VGA_l073_n_151, B1 => VGA_l073_n_150, ZN => VGA_l073_n_161);
  VGA_l073_g12487 : NR3D0BWP7T port map(A1 => VGA_l073_n_148, A2 => VGA_l073_n_87, A3 => VGA_l073_n_40, ZN => VGA_l073_n_160);
  VGA_l073_g12488 : INR2D0BWP7T port map(A1 => VGA_l073_n_44, B1 => VGA_l073_n_149, ZN => VGA_l073_n_159);
  VGA_l073_g12489 : AOI211D0BWP7T port map(A1 => VGA_l073_n_44, A2 => VGA_l073_n_34, B => VGA_l073_n_149, C => VGA_l073_n_98, ZN => VGA_l073_n_158);
  VGA_l073_g12490 : AOI22D0BWP7T port map(A1 => VGA_l073_n_146, A2 => VGA_l073_n_126, B1 => VGA_l073_n_45, B2 => VGA_l073_n_26, ZN => VGA_l073_n_153);
  VGA_l073_g12491 : OAI22D0BWP7T port map(A1 => VGA_l073_n_146, A2 => VGA_l073_n_130, B1 => VGA_l073_n_97, B2 => VGA_x(5), ZN => VGA_l073_n_152);
  VGA_l073_g12492 : INR3D0BWP7T port map(A1 => VGA_l073_n_148, B1 => VGA_l073_n_40, B2 => VGA_l073_n_87, ZN => VGA_l073_n_156);
  VGA_l073_g12493 : AN3D0BWP7T port map(A1 => VGA_l073_n_147, A2 => VGA_l073_n_87, A3 => VGA_l073_n_39, Z => VGA_l073_n_155);
  VGA_l073_g12494 : INR3D0BWP7T port map(A1 => VGA_l073_n_87, B1 => VGA_l073_n_40, B2 => VGA_l073_n_147, ZN => VGA_l073_n_154);
  VGA_l073_g12495 : AN2D1BWP7T port map(A1 => VGA_l073_n_144, A2 => VGA_l073_n_114, Z => VGA_l073_n_151);
  VGA_l073_g12496 : ND2D0BWP7T port map(A1 => VGA_l073_n_143, A2 => VGA_l073_n_113, ZN => VGA_l073_n_150);
  VGA_l073_g12497 : IND4D0BWP7T port map(A1 => VGA_l073_n_108, B1 => VGA_l073_n_109, B2 => VGA_l073_n_106, B3 => VGA_l073_n_107, ZN => VGA_l073_n_149);
  VGA_l073_g12498 : AN3D0BWP7T port map(A1 => VGA_l073_n_128, A2 => VGA_l073_n_70, A3 => VGA_l073_n_76, Z => VGA_l073_n_145);
  VGA_l073_g12499 : OAI221D0BWP7T port map(A1 => VGA_l073_n_101, A2 => y_pos_e3(1), B1 => VGA_l073_n_4, B2 => VGA_l073_n_82, C => VGA_l073_n_100, ZN => VGA_l073_n_148);
  VGA_l073_g12500 : OAI211D0BWP7T port map(A1 => y_pos_e3(1), A2 => VGA_l073_n_41, B => VGA_l073_n_121, C => VGA_l073_n_101, ZN => VGA_l073_n_147);
  VGA_l073_g12501 : MAOI222D0BWP7T port map(A => VGA_x(2), B => x_pos_e3(2), C => VGA_l073_n_83, ZN => VGA_l073_n_146);
  VGA_l073_g12502 : AN3D0BWP7T port map(A1 => VGA_l073_n_124, A2 => VGA_l073_n_94, A3 => VGA_l073_n_92, Z => VGA_l073_n_142);
  VGA_l073_g12503 : INR3D0BWP7T port map(A1 => VGA_l073_n_128, B1 => VGA_l073_n_72, B2 => VGA_l073_n_77, ZN => VGA_l073_n_141);
  VGA_l073_g12504 : AOI211D0BWP7T port map(A1 => VGA_l073_n_101, A2 => VGA_l073_n_100, B => VGA_l073_n_39, C => VGA_l073_n_43, ZN => VGA_l073_n_144);
  VGA_l073_g12505 : AN4D1BWP7T port map(A1 => VGA_l073_n_101, A2 => VGA_l073_n_100, A3 => VGA_l073_n_42, A4 => VGA_l073_n_40, Z => VGA_l073_n_143);
  VGA_l073_g12506 : INR2D0BWP7T port map(A1 => VGA_l073_n_122, B1 => VGA_l073_n_72, ZN => VGA_l073_n_139);
  VGA_l073_g12507 : AN2D1BWP7T port map(A1 => VGA_l073_n_112, A2 => VGA_l073_n_52, Z => VGA_l073_n_138);
  VGA_l073_g12508 : ND2D0BWP7T port map(A1 => VGA_l073_n_123, A2 => VGA_l073_n_131, ZN => VGA_l073_n_137);
  VGA_l073_g12509 : INR2D0BWP7T port map(A1 => VGA_l073_n_104, B1 => VGA_l073_n_1, ZN => VGA_l073_n_140);
  VGA_l073_g12510 : OA221D0BWP7T port map(A1 => VGA_l073_n_67, A2 => VGA_draw_count7(1), B1 => VGA_l073_n_24, B2 => VGA_l073_n_54, C => VGA_l073_n_74, Z => VGA_l073_n_135);
  VGA_l073_g12511 : OAI211D0BWP7T port map(A1 => VGA_draw_count7(1), A2 => VGA_l073_n_58, B => VGA_l073_n_84, C => VGA_l073_n_74, ZN => VGA_l073_n_134);
  VGA_l073_g12512 : OAI211D0BWP7T port map(A1 => VGA_l073_n_13, A2 => VGA_l073_n_54, B => VGA_l073_n_85, C => VGA_l073_n_75, ZN => VGA_l073_n_133);
  VGA_l073_g12513 : OA21D0BWP7T port map(A1 => VGA_l073_n_14, A2 => VGA_l073_n_3, B => VGA_l073_n_124, Z => VGA_l073_n_132);
  VGA_l073_g12514 : ND2D0BWP7T port map(A1 => VGA_l073_n_110, A2 => VGA_l073_n_105, ZN => VGA_l073_n_136);
  VGA_l073_g12515 : CKND1BWP7T port map(I => VGA_l073_n_129, ZN => VGA_l073_n_130);
  VGA_l073_g12516 : CKND1BWP7T port map(I => VGA_l073_n_125, ZN => VGA_l073_n_126);
  VGA_l073_g12517 : IND2D0BWP7T port map(A1 => VGA_l073_n_100, B1 => y_pos_e3(1), ZN => VGA_l073_n_121);
  VGA_l073_g12518 : MOAI22D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l073_n_10, B1 => VGA_l073_n_49, B2 => VGA_l073_n_32, ZN => VGA_l073_n_120);
  VGA_l073_g12519 : AOI21D0BWP7T port map(A1 => VGA_l073_n_59, A2 => VGA_l073_n_27, B => VGA_l073_n_93, ZN => VGA_l073_n_119);
  VGA_l073_g12520 : AOI211D0BWP7T port map(A1 => VGA_l073_n_55, A2 => VGA_l073_n_24, B => VGA_l073_n_93, C => VGA_l073_n_78, ZN => VGA_l073_n_118);
  VGA_l073_g12521 : OAI221D0BWP7T port map(A1 => VGA_l073_n_62, A2 => VGA_l073_n_0, B1 => VGA_l073_n_29, B2 => VGA_l073_n_64, C => VGA_l073_n_92, ZN => VGA_l073_n_117);
  VGA_l073_g12522 : OA21D0BWP7T port map(A1 => VGA_l073_n_62, A2 => VGA_l073_n_64, B => VGA_l073_n_92, Z => VGA_l073_n_131);
  VGA_l073_g12523 : AOI22D0BWP7T port map(A1 => VGA_l073_n_66, A2 => VGA_l073_n_31, B1 => VGA_l073_n_47, B2 => VGA_x(2), ZN => VGA_l073_n_129);
  VGA_l073_g12524 : NR3D0BWP7T port map(A1 => VGA_l073_n_80, A2 => VGA_l073_n_73, A3 => VGA_l073_n_61, ZN => VGA_l073_n_128);
  VGA_l073_g12525 : IND2D0BWP7T port map(A1 => VGA_l073_n_37, B1 => VGA_l073_n_102, ZN => VGA_l073_n_127);
  VGA_l073_g12526 : OAI22D0BWP7T port map(A1 => VGA_l073_n_66, A2 => VGA_l073_n_31, B1 => VGA_l073_n_47, B2 => VGA_x(2), ZN => VGA_l073_n_125);
  VGA_l073_g12527 : AN3D0BWP7T port map(A1 => VGA_l073_n_68, A2 => VGA_l073_n_75, A3 => VGA_l073_n_69, Z => VGA_l073_n_124);
  VGA_l073_g12528 : AN2D1BWP7T port map(A1 => VGA_l073_n_88, A2 => VGA_l073_n_68, Z => VGA_l073_n_123);
  VGA_l073_g12529 : AN2D1BWP7T port map(A1 => VGA_l073_n_89, A2 => VGA_l073_n_58, Z => VGA_l073_n_122);
  VGA_l073_g12530 : AOI221D0BWP7T port map(A1 => VGA_l073_n_61, A2 => VGA_draw_count7(0), B1 => VGA_l073_n_56, B2 => VGA_l073_n_25, C => VGA_l073_n_80, ZN => VGA_l073_n_112);
  VGA_l073_g12531 : AO222D0BWP7T port map(A1 => VGA_l073_n_61, A2 => VGA_l073_n_24, B1 => VGA_l073_n_55, B2 => VGA_l073_n_13, C1 => VGA_l073_n_53, C2 => VGA_l073_n_27, Z => VGA_l073_n_111);
  VGA_l073_g12532 : OAI22D0BWP7T port map(A1 => VGA_l073_n_45, A2 => VGA_l073_n_26, B1 => VGA_l073_n_46, B2 => VGA_l073_n_16, ZN => VGA_l073_n_110);
  VGA_l073_g12533 : MAOI22D0BWP7T port map(A1 => VGA_l073_n_50, A2 => VGA_l073_n_35, B1 => VGA_l073_n_50, B2 => VGA_l073_n_35, ZN => VGA_l073_n_109);
  VGA_l073_g12534 : OAI22D0BWP7T port map(A1 => VGA_l073_n_65, A2 => VGA_l073_n_15, B1 => VGA_l073_n_36, B2 => VGA_y(9), ZN => VGA_l073_n_108);
  VGA_l073_g12535 : AOI22D0BWP7T port map(A1 => VGA_l073_n_65, A2 => VGA_l073_n_15, B1 => VGA_l073_n_36, B2 => VGA_y(9), ZN => VGA_l073_n_107);
  VGA_l073_g12536 : MAOI22D0BWP7T port map(A1 => VGA_l073_n_48, A2 => VGA_l073_n_28, B1 => VGA_l073_n_48, B2 => VGA_l073_n_28, ZN => VGA_l073_n_106);
  VGA_l073_g12538 : MAOI22D0BWP7T port map(A1 => VGA_l073_n_38, A2 => VGA_l073_n_19, B1 => VGA_l073_n_38, B2 => VGA_l073_n_19, ZN => VGA_l073_n_116);
  VGA_l073_g12540 : MOAI22D0BWP7T port map(A1 => VGA_l073_n_38, A2 => VGA_l073_n_22, B1 => VGA_l073_n_38, B2 => VGA_l073_n_22, ZN => VGA_l073_n_115);
  VGA_l073_g12541 : MAOI22D0BWP7T port map(A1 => VGA_l073_n_37, A2 => VGA_l073_n_33, B1 => VGA_l073_n_37, B2 => VGA_l073_n_33, ZN => VGA_l073_n_114);
  VGA_l073_g12542 : MOAI22D0BWP7T port map(A1 => VGA_l073_n_37, A2 => VGA_l073_n_23, B1 => VGA_l073_n_37, B2 => VGA_l073_n_23, ZN => VGA_l073_n_113);
  VGA_l073_g12543 : AOI21D0BWP7T port map(A1 => VGA_l073_n_56, A2 => VGA_l073_n_24, B => VGA_l073_n_63, ZN => VGA_l073_n_99);
  VGA_l073_g12544 : NR2D0BWP7T port map(A1 => VGA_l073_n_44, A2 => VGA_l073_n_34, ZN => VGA_l073_n_98);
  VGA_l073_g12545 : IND2D0BWP7T port map(A1 => VGA_l073_n_46, B1 => x_pos_e3(5), ZN => VGA_l073_n_97);
  VGA_l073_g12546 : ND2D0BWP7T port map(A1 => VGA_l073_n_46, A2 => VGA_l073_n_16, ZN => VGA_l073_n_105);
  VGA_l073_g12547 : NR2D0BWP7T port map(A1 => VGA_l073_n_66, A2 => VGA_l073_n_31, ZN => VGA_l073_n_96);
  VGA_l073_g12548 : NR2D0BWP7T port map(A1 => VGA_l073_n_71, A2 => VGA_l073_n_41, ZN => VGA_l073_n_104);
  VGA_l073_g12550 : NR2D0BWP7T port map(A1 => VGA_l073_n_79, A2 => VGA_l073_n_78, ZN => VGA_l073_n_103);
  VGA_l073_g12551 : NR2D0BWP7T port map(A1 => VGA_l073_n_71, A2 => VGA_l073_n_82, ZN => VGA_l073_n_102);
  VGA_l073_g12552 : ND2D0BWP7T port map(A1 => VGA_l073_n_82, A2 => VGA_y(1), ZN => VGA_l073_n_101);
  VGA_l073_g12553 : IND2D0BWP7T port map(A1 => VGA_y(1), B1 => VGA_l073_n_41, ZN => VGA_l073_n_100);
  VGA_l073_g12554 : CKND1BWP7T port map(I => VGA_l073_n_90, ZN => VGA_l073_n_91);
  VGA_l073_g12555 : AOI21D0BWP7T port map(A1 => VGA_l073_n_59, A2 => VGA_l073_n_25, B => VGA_l073_n_73, ZN => VGA_l073_n_86);
  VGA_l073_g12556 : OAI21D0BWP7T port map(A1 => VGA_l073_n_56, A2 => VGA_l073_n_53, B => VGA_l073_n_24, ZN => VGA_l073_n_85);
  VGA_l073_g12557 : AO21D0BWP7T port map(A1 => VGA_l073_n_60, A2 => VGA_l073_n_54, B => VGA_l073_n_62, Z => VGA_l073_n_84);
  VGA_l073_g12558 : IAO21D0BWP7T port map(A1 => VGA_l073_n_60, A2 => VGA_l073_n_13, B => VGA_l073_n_55, ZN => VGA_l073_n_94);
  VGA_l073_g12559 : OAI21D0BWP7T port map(A1 => VGA_l073_n_52, A2 => VGA_draw_count7(1), B => VGA_l073_n_70, ZN => VGA_l073_n_93);
  VGA_l073_g12560 : AOI22D0BWP7T port map(A1 => VGA_l073_n_51, A2 => VGA_x(0), B1 => VGA_x(1), B2 => VGA_l073_n_6, ZN => VGA_l073_n_83);
  VGA_l073_g12561 : OA22D0BWP7T port map(A1 => VGA_l073_n_64, A2 => VGA_l073_n_12, B1 => VGA_l073_n_25, B2 => VGA_l073_n_0, Z => VGA_l073_n_92);
  VGA_l073_g12562 : OAI21D0BWP7T port map(A1 => VGA_l073_n_57, A2 => VGA_l073_n_13, B => VGA_l073_n_69, ZN => VGA_l073_n_90);
  VGA_l073_g12563 : AOI22D0BWP7T port map(A1 => VGA_l073_n_56, A2 => VGA_l073_n_13, B1 => VGA_l073_n_59, B2 => VGA_l073_n_24, ZN => VGA_l073_n_89);
  VGA_l073_g12564 : IAO21D0BWP7T port map(A1 => VGA_l073_n_0, A2 => VGA_l073_n_24, B => VGA_l073_n_79, ZN => VGA_l073_n_88);
  VGA_l073_g12565 : MOAI22D0BWP7T port map(A1 => VGA_l073_n_43, A2 => VGA_y(0), B1 => VGA_l073_n_43, B2 => VGA_y(0), ZN => VGA_l073_n_87);
  VGA_l073_g12568 : INVD0BWP7T port map(I => VGA_l073_n_41, ZN => VGA_l073_n_82);
  VGA_l073_g12569 : CKND1BWP7T port map(I => VGA_l073_n_26, ZN => VGA_l073_n_81);
  VGA_l073_g12570 : NR2D0BWP7T port map(A1 => VGA_l073_n_54, A2 => VGA_draw_count7(1), ZN => VGA_l073_n_80);
  VGA_l073_g12571 : INR2D0BWP7T port map(A1 => VGA_l073_n_63, B1 => VGA_l073_n_25, ZN => VGA_l073_n_79);
  VGA_l073_g12572 : NR2D0BWP7T port map(A1 => VGA_l073_n_0, A2 => VGA_draw_count7(1), ZN => VGA_l073_n_78);
  VGA_l073_g12573 : NR2D0BWP7T port map(A1 => VGA_l073_n_57, A2 => VGA_l073_n_29, ZN => VGA_l073_n_77);
  VGA_l073_g12574 : ND2D0BWP7T port map(A1 => VGA_l073_n_55, A2 => VGA_draw_count7(1), ZN => VGA_l073_n_76);
  VGA_l073_g12575 : ND2D0BWP7T port map(A1 => VGA_l073_n_53, A2 => VGA_l073_n_13, ZN => VGA_l073_n_75);
  VGA_l073_g12576 : ND2D0BWP7T port map(A1 => VGA_l073_n_53, A2 => VGA_draw_count7(1), ZN => VGA_l073_n_74);
  VGA_l073_g12577 : NR2D0BWP7T port map(A1 => VGA_l073_n_56, A2 => VGA_l073_n_59, ZN => VGA_l073_n_67);
  VGA_l073_g12578 : AN2D1BWP7T port map(A1 => VGA_l073_n_63, A2 => VGA_l073_n_27, Z => VGA_l073_n_73);
  VGA_l073_g12579 : NR2D0BWP7T port map(A1 => VGA_l073_n_52, A2 => VGA_l073_n_13, ZN => VGA_l073_n_72);
  VGA_l073_g12580 : ND2D0BWP7T port map(A1 => VGA_l073_n_40, A2 => VGA_l073_n_43, ZN => VGA_l073_n_71);
  VGA_l073_g12581 : IND2D0BWP7T port map(A1 => VGA_l073_n_62, B1 => VGA_l073_n_56, ZN => VGA_l073_n_70);
  VGA_l073_g12582 : ND2D0BWP7T port map(A1 => VGA_l073_n_63, A2 => VGA_l073_n_13, ZN => VGA_l073_n_69);
  VGA_l073_g12583 : IND2D0BWP7T port map(A1 => VGA_l073_n_62, B1 => VGA_l073_n_63, ZN => VGA_l073_n_68);
  VGA_l073_g12584 : INVD0BWP7T port map(I => VGA_l073_n_61, ZN => VGA_l073_n_60);
  VGA_l073_g12585 : INVD0BWP7T port map(I => VGA_l073_n_59, ZN => VGA_l073_n_58);
  VGA_l073_g12586 : INVD1BWP7T port map(I => VGA_l073_n_57, ZN => VGA_l073_n_56);
  VGA_l073_g12587 : INVD0BWP7T port map(I => VGA_l073_n_55, ZN => VGA_l073_n_54);
  VGA_l073_g12588 : INVD0BWP7T port map(I => VGA_l073_n_53, ZN => VGA_l073_n_52);
  VGA_l073_g12589 : IAO21D0BWP7T port map(A1 => VGA_x(1), A2 => VGA_l073_n_6, B => x_pos_e3(0), ZN => VGA_l073_n_51);
  VGA_l073_g12590 : OAI21D0BWP7T port map(A1 => VGA_l073_n_7, A2 => x_pos_e3(4), B => VGA_l073_n_26, ZN => VGA_l073_n_66);
  VGA_l073_g12591 : AOI21D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l073_n_5, B => VGA_l073_n_28, ZN => VGA_l073_n_65);
  VGA_l073_g12592 : IND2D0BWP7T port map(A1 => VGA_l073_n_30, B1 => VGA_draw_count7(4), ZN => VGA_l073_n_64);
  VGA_l073_g12593 : INR2D0BWP7T port map(A1 => VGA_draw_count7(4), B1 => VGA_l073_n_17, ZN => VGA_l073_n_63);
  VGA_l073_g12594 : INR2D0BWP7T port map(A1 => VGA_l073_n_29, B1 => VGA_l073_n_27, ZN => VGA_l073_n_62);
  VGA_l073_g12596 : NR2D0BWP7T port map(A1 => VGA_l073_n_14, A2 => VGA_draw_count7(4), ZN => VGA_l073_n_61);
  VGA_l073_g12597 : NR2D0BWP7T port map(A1 => VGA_l073_n_30, A2 => VGA_draw_count7(4), ZN => VGA_l073_n_59);
  VGA_l073_g12598 : IND2D0BWP7T port map(A1 => VGA_l073_n_14, B1 => VGA_draw_count7(4), ZN => VGA_l073_n_57);
  VGA_l073_g12599 : NR2D0BWP7T port map(A1 => VGA_l073_n_17, A2 => VGA_draw_count7(4), ZN => VGA_l073_n_55);
  VGA_l073_g12600 : NR2D0BWP7T port map(A1 => VGA_l073_n_18, A2 => VGA_draw_count7(4), ZN => VGA_l073_n_53);
  VGA_l073_g12601 : CKND1BWP7T port map(I => VGA_l073_n_43, ZN => VGA_l073_n_42);
  VGA_l073_g12602 : CKND1BWP7T port map(I => VGA_l073_n_40, ZN => VGA_l073_n_39);
  VGA_l073_g12603 : MOAI22D0BWP7T port map(A1 => VGA_y(8), A2 => y_pos_e3(8), B1 => VGA_y(8), B2 => y_pos_e3(8), ZN => VGA_l073_n_50);
  VGA_l073_g12604 : MOAI22D0BWP7T port map(A1 => VGA_x(7), A2 => x_pos_e3(7), B1 => VGA_x(7), B2 => x_pos_e3(7), ZN => VGA_l073_n_49);
  VGA_l073_g12605 : MOAI22D0BWP7T port map(A1 => VGA_y(7), A2 => y_pos_e3(7), B1 => VGA_y(7), B2 => y_pos_e3(7), ZN => VGA_l073_n_48);
  VGA_l073_g12606 : MAOI22D0BWP7T port map(A1 => VGA_x(3), A2 => x_pos_e3(3), B1 => VGA_x(3), B2 => x_pos_e3(3), ZN => VGA_l073_n_47);
  VGA_l073_g12607 : MOAI22D0BWP7T port map(A1 => VGA_x(6), A2 => x_pos_e3(6), B1 => VGA_x(6), B2 => x_pos_e3(6), ZN => VGA_l073_n_46);
  VGA_l073_g12608 : MOAI22D0BWP7T port map(A1 => VGA_x(5), A2 => x_pos_e3(5), B1 => VGA_x(5), B2 => x_pos_e3(5), ZN => VGA_l073_n_45);
  VGA_l073_g12609 : MAOI22D0BWP7T port map(A1 => VGA_y(5), A2 => y_pos_e3(5), B1 => VGA_y(5), B2 => y_pos_e3(5), ZN => VGA_l073_n_44);
  VGA_l073_g12610 : MOAI22D0BWP7T port map(A1 => VGA_y(1), A2 => y_pos_e3(1), B1 => VGA_y(1), B2 => y_pos_e3(1), ZN => VGA_l073_n_43);
  VGA_l073_g12611 : MOAI22D0BWP7T port map(A1 => VGA_y(2), A2 => y_pos_e3(2), B1 => VGA_y(2), B2 => y_pos_e3(2), ZN => VGA_l073_n_41);
  VGA_l073_g12612 : MOAI22D0BWP7T port map(A1 => VGA_y(0), A2 => y_pos_e3(0), B1 => VGA_y(0), B2 => y_pos_e3(0), ZN => VGA_l073_n_40);
  VGA_l073_g12613 : MAOI22D0BWP7T port map(A1 => VGA_y(4), A2 => y_pos_e3(4), B1 => VGA_y(4), B2 => y_pos_e3(4), ZN => VGA_l073_n_38);
  VGA_l073_g12614 : MOAI22D0BWP7T port map(A1 => VGA_y(3), A2 => y_pos_e3(3), B1 => VGA_y(3), B2 => y_pos_e3(3), ZN => VGA_l073_n_37);
  VGA_l073_g12615 : INVD1BWP7T port map(I => VGA_l073_n_25, ZN => VGA_l073_n_24);
  VGA_l073_g12616 : IND2D0BWP7T port map(A1 => VGA_y(8), B1 => y_pos_e3(8), ZN => VGA_l073_n_36);
  VGA_l073_g12617 : INR2D0BWP7T port map(A1 => y_pos_e3(7), B1 => VGA_y(7), ZN => VGA_l073_n_35);
  VGA_l073_g12618 : IND2D0BWP7T port map(A1 => y_pos_e3(4), B1 => VGA_y(4), ZN => VGA_l073_n_34);
  VGA_l073_g12619 : IND2D0BWP7T port map(A1 => y_pos_e3(2), B1 => VGA_y(2), ZN => VGA_l073_n_33);
  VGA_l073_g12620 : IND2D0BWP7T port map(A1 => x_pos_e3(6), B1 => VGA_x(6), ZN => VGA_l073_n_32);
  VGA_l073_g12621 : IND2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_e3(3), ZN => VGA_l073_n_31);
  VGA_l073_g12622 : ND2D0BWP7T port map(A1 => VGA_draw_count7(2), A2 => VGA_draw_count7(3), ZN => VGA_l073_n_30);
  VGA_l073_g12623 : ND2D0BWP7T port map(A1 => VGA_l073_n_3, A2 => VGA_draw_count7(0), ZN => VGA_l073_n_29);
  VGA_l073_g12624 : NR2D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l073_n_5, ZN => VGA_l073_n_28);
  VGA_l073_g12625 : NR2D0BWP7T port map(A1 => VGA_l073_n_3, A2 => VGA_draw_count7(0), ZN => VGA_l073_n_27);
  VGA_l073_g12626 : ND2D0BWP7T port map(A1 => VGA_l073_n_7, A2 => x_pos_e3(4), ZN => VGA_l073_n_26);
  VGA_l073_g12627 : ND2D0BWP7T port map(A1 => VGA_draw_count7(1), A2 => VGA_draw_count7(0), ZN => VGA_l073_n_25);
  VGA_l073_g12629 : CKND1BWP7T port map(I => VGA_l073_n_13, ZN => VGA_l073_n_12);
  VGA_l073_g12630 : IND2D0BWP7T port map(A1 => VGA_y(4), B1 => y_pos_e3(4), ZN => VGA_l073_n_11);
  VGA_l073_g12631 : ND2D0BWP7T port map(A1 => VGA_l073_n_8, A2 => y_pos_e3(2), ZN => VGA_l073_n_23);
  VGA_l073_g12632 : NR2D0BWP7T port map(A1 => VGA_l073_n_9, A2 => y_pos_e3(3), ZN => VGA_l073_n_22);
  VGA_l073_g12633 : INR2D0BWP7T port map(A1 => x_pos_e3(7), B1 => VGA_x(7), ZN => VGA_l073_n_21);
  VGA_l073_g12634 : ND2D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l073_n_10, ZN => VGA_l073_n_20);
  VGA_l073_g12635 : INR2D0BWP7T port map(A1 => y_pos_e3(3), B1 => VGA_y(3), ZN => VGA_l073_n_19);
  VGA_l073_g12636 : IND2D0BWP7T port map(A1 => VGA_draw_count7(2), B1 => VGA_draw_count7(3), ZN => VGA_l073_n_18);
  VGA_l073_g12637 : IND2D0BWP7T port map(A1 => VGA_draw_count7(3), B1 => VGA_draw_count7(2), ZN => VGA_l073_n_17);
  VGA_l073_g12638 : INR2D0BWP7T port map(A1 => VGA_x(5), B1 => x_pos_e3(5), ZN => VGA_l073_n_16);
  VGA_l073_g12639 : IND2D0BWP7T port map(A1 => y_pos_e3(5), B1 => VGA_y(5), ZN => VGA_l073_n_15);
  VGA_l073_g12640 : OR2D0BWP7T port map(A1 => VGA_draw_count7(2), A2 => VGA_draw_count7(3), Z => VGA_l073_n_14);
  VGA_l073_g12641 : NR2D0BWP7T port map(A1 => VGA_draw_count7(1), A2 => VGA_draw_count7(0), ZN => VGA_l073_n_13);
  VGA_l073_g12642 : CKND1BWP7T port map(I => x_pos_e3(8), ZN => VGA_l073_n_10);
  VGA_l073_g12643 : CKND1BWP7T port map(I => VGA_y(3), ZN => VGA_l073_n_9);
  VGA_l073_g12644 : CKND1BWP7T port map(I => VGA_y(2), ZN => VGA_l073_n_8);
  VGA_l073_g12645 : CKND1BWP7T port map(I => VGA_x(4), ZN => VGA_l073_n_7);
  VGA_l073_g12646 : CKND1BWP7T port map(I => x_pos_e3(1), ZN => VGA_l073_n_6);
  VGA_l073_g12647 : CKND1BWP7T port map(I => y_pos_e3(6), ZN => VGA_l073_n_5);
  VGA_l073_g12648 : CKND1BWP7T port map(I => y_pos_e3(1), ZN => VGA_l073_n_4);
  VGA_l073_g12649 : INVD0BWP7T port map(I => VGA_draw_count7(1), ZN => VGA_l073_n_3);
  VGA_l073_g2 : MUX2ND0BWP7T port map(I0 => VGA_y(3), I1 => VGA_l073_n_9, S => VGA_l073_n_38, ZN => VGA_l073_n_2);
  VGA_l073_g12650 : MUX2ND0BWP7T port map(I0 => VGA_l073_n_8, I1 => VGA_y(2), S => VGA_l073_n_37, ZN => VGA_l073_n_1);
  VGA_l073_g12651 : IND2D1BWP7T port map(A1 => VGA_l073_n_18, B1 => VGA_draw_count7(4), ZN => VGA_l073_n_0);
  VGA_l073_g12652 : INVD0BWP7T port map(I => VGA_l073_n_66, ZN => VGA_l073_n_95);
  VGA_l074_g12402 : OAI211D0BWP7T port map(A1 => VGA_l074_n_76, A2 => VGA_l074_n_195, B => VGA_l074_n_243, C => VGA_l074_n_223, ZN => VGA_r8);
  VGA_l074_g12403 : AOI211D0BWP7T port map(A1 => VGA_l074_n_206, A2 => VGA_l074_n_111, B => VGA_l074_n_242, C => VGA_l074_n_225, ZN => VGA_l074_n_243);
  VGA_l074_g12404 : OAI211D0BWP7T port map(A1 => VGA_l074_n_162, A2 => VGA_l074_n_216, B => VGA_l074_n_241, C => VGA_l074_n_238, ZN => VGA_l074_n_242);
  VGA_l074_g12405 : NR4D0BWP7T port map(A1 => VGA_l074_n_239, A2 => VGA_l074_n_227, A3 => VGA_l074_n_219, A4 => VGA_l074_n_220, ZN => VGA_l074_n_241);
  VGA_l074_g12406 : OAI211D0BWP7T port map(A1 => VGA_l074_n_91, A2 => VGA_l074_n_212, B => VGA_l074_n_237, C => VGA_l074_n_235, ZN => VGA_g8);
  VGA_l074_g12407 : NR4D0BWP7T port map(A1 => VGA_l074_n_233, A2 => VGA_l074_n_191, A3 => VGA_l074_n_151, A4 => VGA_l074_n_138, ZN => VGA_l074_n_239);
  VGA_l074_g12408 : NR4D0BWP7T port map(A1 => VGA_l074_n_226, A2 => VGA_l074_n_228, A3 => VGA_l074_n_221, A4 => VGA_l074_n_192, ZN => VGA_l074_n_238);
  VGA_l074_g12409 : AOI211D0BWP7T port map(A1 => VGA_l074_n_206, A2 => VGA_l074_n_117, B => VGA_l074_n_236, C => VGA_l074_n_218, ZN => VGA_l074_n_237);
  VGA_l074_g12410 : OAI211D0BWP7T port map(A1 => VGA_l074_n_99, A2 => VGA_l074_n_195, B => VGA_l074_n_230, C => VGA_l074_n_224, ZN => VGA_l074_n_236);
  VGA_l074_g12411 : AOI211D0BWP7T port map(A1 => VGA_l074_n_211, A2 => VGA_l074_n_137, B => VGA_l074_n_231, C => VGA_l074_n_213, ZN => VGA_l074_n_235);
  VGA_l074_g12412 : OAI32D0BWP7T port map(A1 => VGA_l074_n_24, A2 => VGA_l074_n_60, A3 => VGA_l074_n_216, B1 => VGA_l074_n_94, B2 => VGA_l074_n_215, ZN => VGA_b8);
  VGA_l074_g12413 : ND4D0BWP7T port map(A1 => VGA_l074_n_210, A2 => VGA_l074_n_189, A3 => VGA_l074_n_176, A4 => VGA_l074_n_165, ZN => VGA_l074_n_233);
  VGA_l074_g12414 : OAI211D0BWP7T port map(A1 => VGA_l074_n_191, A2 => VGA_l074_n_209, B => VGA_l074_n_204, C => VGA_l074_n_199, ZN => VGA_enable8);
  VGA_l074_g12415 : OAI22D0BWP7T port map(A1 => VGA_l074_n_217, A2 => VGA_l074_n_139, B1 => VGA_l074_n_207, B2 => VGA_l074_n_131, ZN => VGA_l074_n_231);
  VGA_l074_g12416 : AOI31D0BWP7T port map(A1 => VGA_l074_n_190, A2 => VGA_l074_n_182, A3 => VGA_l074_n_77, B => VGA_l074_n_229, ZN => VGA_l074_n_230);
  VGA_l074_g12417 : AOI21D0BWP7T port map(A1 => VGA_l074_n_103, A2 => VGA_l074_n_86, B => VGA_l074_n_216, ZN => VGA_l074_n_229);
  VGA_l074_g12418 : AOI31D0BWP7T port map(A1 => VGA_l074_n_145, A2 => VGA_l074_n_88, A3 => VGA_l074_n_75, B => VGA_l074_n_217, ZN => VGA_l074_n_228);
  VGA_l074_g12419 : AOI31D0BWP7T port map(A1 => VGA_l074_n_122, A2 => VGA_l074_n_118, A3 => VGA_l074_n_60, B => VGA_l074_n_214, ZN => VGA_l074_n_227);
  VGA_l074_g12420 : AOI31D0BWP7T port map(A1 => VGA_l074_n_142, A2 => VGA_l074_n_122, A3 => VGA_l074_n_88, B => VGA_l074_n_215, ZN => VGA_l074_n_226);
  VGA_l074_g12421 : AOI22D0BWP7T port map(A1 => VGA_l074_n_205, A2 => VGA_l074_n_195, B1 => VGA_l074_n_119, B2 => VGA_l074_n_89, ZN => VGA_l074_n_225);
  VGA_l074_g12422 : AO21D0BWP7T port map(A1 => VGA_l074_n_123, A2 => VGA_l074_n_91, B => VGA_l074_n_215, Z => VGA_l074_n_224);
  VGA_l074_g12423 : OA21D0BWP7T port map(A1 => VGA_l074_n_208, A2 => VGA_l074_n_157, B => VGA_l074_n_222, Z => VGA_l074_n_223);
  VGA_l074_g12424 : AO31D0BWP7T port map(A1 => VGA_l074_n_135, A2 => VGA_l074_n_68, A3 => VGA_l074_n_69, B => VGA_l074_n_204, Z => VGA_l074_n_222);
  VGA_l074_g12425 : AOI21D0BWP7T port map(A1 => VGA_l074_n_89, A2 => VGA_l074_n_52, B => VGA_l074_n_212, ZN => VGA_l074_n_221);
  VGA_l074_g12426 : AOI31D0BWP7T port map(A1 => VGA_l074_n_132, A2 => VGA_l074_n_76, A3 => VGA_l074_n_58, B => VGA_l074_n_207, ZN => VGA_l074_n_220);
  VGA_l074_g12427 : OA21D0BWP7T port map(A1 => VGA_l074_n_134, A2 => VGA_l074_n_90, B => VGA_l074_n_211, Z => VGA_l074_n_219);
  VGA_l074_g12428 : AOI21D0BWP7T port map(A1 => VGA_l074_n_88, A2 => VGA_l074_n_0, B => VGA_l074_n_204, ZN => VGA_l074_n_218);
  VGA_l074_g12429 : AOI32D0BWP7T port map(A1 => VGA_l074_n_190, A2 => VGA_l074_n_181, A3 => VGA_l074_n_38, B1 => VGA_l074_n_202, B2 => VGA_l074_n_154, ZN => VGA_l074_n_214);
  VGA_l074_g12430 : AOI21D0BWP7T port map(A1 => VGA_l074_n_103, A2 => VGA_l074_n_68, B => VGA_l074_n_208, ZN => VGA_l074_n_213);
  VGA_l074_g12431 : AOI22D0BWP7T port map(A1 => VGA_l074_n_203, A2 => VGA_l074_n_156, B1 => VGA_l074_n_202, B2 => VGA_l074_n_143, ZN => VGA_l074_n_217);
  VGA_l074_g12432 : AOI22D0BWP7T port map(A1 => VGA_l074_n_202, A2 => VGA_l074_n_160, B1 => VGA_l074_n_203, B2 => VGA_l074_n_144, ZN => VGA_l074_n_216);
  VGA_l074_g12433 : AOI32D0BWP7T port map(A1 => VGA_l074_n_198, A2 => VGA_l074_n_1, A3 => VGA_l074_n_104, B1 => VGA_l074_n_203, B2 => VGA_l074_n_155, ZN => VGA_l074_n_215);
  VGA_l074_g12434 : OAI31D0BWP7T port map(A1 => VGA_l074_n_2, A2 => VGA_l074_n_127, A3 => VGA_l074_n_179, B => VGA_l074_n_201, ZN => VGA_l074_n_210);
  VGA_l074_g12435 : NR4D0BWP7T port map(A1 => VGA_l074_n_200, A2 => VGA_l074_n_186, A3 => VGA_l074_n_182, A4 => VGA_l074_n_185, ZN => VGA_l074_n_209);
  VGA_l074_g12436 : MAOI22D0BWP7T port map(A1 => VGA_l074_n_196, A2 => VGA_l074_n_170, B1 => VGA_l074_n_191, B2 => VGA_l074_n_165, ZN => VGA_l074_n_212);
  VGA_l074_g12437 : OAI22D0BWP7T port map(A1 => VGA_l074_n_197, A2 => VGA_l074_n_171, B1 => VGA_l074_n_193, B2 => VGA_l074_n_150, ZN => VGA_l074_n_211);
  VGA_l074_g12438 : CKND1BWP7T port map(I => VGA_l074_n_206, ZN => VGA_l074_n_205);
  VGA_l074_g12439 : AOI22D0BWP7T port map(A1 => VGA_l074_n_196, A2 => VGA_l074_n_169, B1 => VGA_l074_n_194, B2 => VGA_l074_n_151, ZN => VGA_l074_n_208);
  VGA_l074_g12440 : MAOI22D0BWP7T port map(A1 => VGA_l074_n_196, A2 => VGA_l074_n_151, B1 => VGA_l074_n_193, B2 => VGA_l074_n_168, ZN => VGA_l074_n_207);
  VGA_l074_g12441 : OAI22D0BWP7T port map(A1 => VGA_l074_n_197, A2 => VGA_l074_n_167, B1 => VGA_l074_n_191, B2 => VGA_l074_n_176, ZN => VGA_l074_n_206);
  VGA_l074_g12442 : MAOI22D0BWP7T port map(A1 => VGA_l074_n_196, A2 => VGA_l074_n_140, B1 => VGA_l074_n_193, B2 => VGA_l074_n_167, ZN => VGA_l074_n_204);
  VGA_l074_g12443 : INR2D0BWP7T port map(A1 => VGA_l074_n_198, B1 => VGA_l074_n_114, ZN => VGA_l074_n_203);
  VGA_l074_g12444 : INR2D0BWP7T port map(A1 => VGA_l074_n_198, B1 => VGA_l074_n_113, ZN => VGA_l074_n_202);
  VGA_l074_g12445 : CKND1BWP7T port map(I => VGA_l074_n_200, ZN => VGA_l074_n_201);
  VGA_l074_g12446 : OAI21D0BWP7T port map(A1 => VGA_l074_n_177, A2 => VGA_l074_n_161, B => VGA_l074_n_194, ZN => VGA_l074_n_199);
  VGA_l074_g12447 : ND3D0BWP7T port map(A1 => VGA_l074_n_188, A2 => VGA_l074_n_176, A3 => VGA_l074_n_165, ZN => VGA_l074_n_200);
  VGA_l074_g12448 : INVD0BWP7T port map(I => VGA_l074_n_197, ZN => VGA_l074_n_196);
  VGA_l074_g12449 : INR2D0BWP7T port map(A1 => VGA_l074_n_185, B1 => VGA_l074_n_191, ZN => VGA_l074_n_198);
  VGA_l074_g12450 : ND2D0BWP7T port map(A1 => VGA_l074_n_190, A2 => VGA_l074_n_184, ZN => VGA_l074_n_197);
  VGA_l074_g12451 : CKND1BWP7T port map(I => VGA_l074_n_193, ZN => VGA_l074_n_194);
  VGA_l074_g12452 : AOI211D0BWP7T port map(A1 => VGA_l074_n_122, A2 => VGA_l074_n_74, B => VGA_l074_n_191, C => VGA_l074_n_183, ZN => VGA_l074_n_192);
  VGA_l074_g12453 : IND2D0BWP7T port map(A1 => VGA_l074_n_189, B1 => VGA_l074_n_190, ZN => VGA_l074_n_195);
  VGA_l074_g12454 : ND2D0BWP7T port map(A1 => VGA_l074_n_190, A2 => VGA_l074_n_164, ZN => VGA_l074_n_193);
  VGA_l074_g12455 : INVD1BWP7T port map(I => VGA_l074_n_191, ZN => VGA_l074_n_190);
  VGA_l074_g12456 : OAI221D0BWP7T port map(A1 => VGA_l074_n_49, A2 => VGA_l074_n_32, B1 => VGA_l074_n_20, B2 => VGA_l074_n_21, C => VGA_l074_n_187, ZN => VGA_l074_n_191);
  VGA_l074_g12457 : AOI22D0BWP7T port map(A1 => VGA_l074_n_184, A2 => VGA_l074_n_161, B1 => VGA_l074_n_170, B2 => VGA_l074_n_164, ZN => VGA_l074_n_188);
  VGA_l074_g12458 : AOI33D0BWP7T port map(A1 => VGA_l074_n_184, A2 => VGA_l074_n_143, A3 => VGA_l074_n_113, B1 => VGA_l074_n_164, B2 => VGA_l074_n_156, B3 => VGA_l074_n_114, ZN => VGA_l074_n_189);
  VGA_l074_g12459 : AOI211D0BWP7T port map(A1 => VGA_l074_n_173, A2 => VGA_l074_n_136, B => VGA_l074_n_178, C => VGA_l074_n_120, ZN => VGA_l074_n_187);
  VGA_l074_g12460 : OA21D0BWP7T port map(A1 => VGA_l074_n_180, A2 => VGA_l074_n_170, B => VGA_l074_n_184, Z => VGA_l074_n_186);
  VGA_l074_g12461 : NR2D0BWP7T port map(A1 => VGA_l074_n_179, A2 => VGA_l074_n_115, ZN => VGA_l074_n_185);
  VGA_l074_g12462 : NR2D0BWP7T port map(A1 => VGA_l074_n_179, A2 => VGA_l074_n_116, ZN => VGA_l074_n_184);
  VGA_l074_g12463 : CKND1BWP7T port map(I => VGA_l074_n_182, ZN => VGA_l074_n_183);
  VGA_l074_g12464 : AO32D0BWP7T port map(A1 => VGA_l074_n_166, A2 => VGA_l074_n_102, A3 => VGA_l074_n_37, B1 => VGA_l074_n_175, B2 => VGA_y(4), Z => VGA_l074_n_181);
  VGA_l074_g12465 : OAI22D0BWP7T port map(A1 => VGA_l074_n_172, A2 => VGA_l074_n_113, B1 => VGA_l074_n_174, B2 => VGA_l074_n_38, ZN => VGA_l074_n_182);
  VGA_l074_g12466 : IND2D0BWP7T port map(A1 => VGA_l074_n_177, B1 => VGA_l074_n_167, ZN => VGA_l074_n_180);
  VGA_l074_g12467 : MOAI22D0BWP7T port map(A1 => VGA_l074_n_163, A2 => VGA_l074_n_136, B1 => VGA_l074_n_21, B2 => VGA_l074_n_20, ZN => VGA_l074_n_178);
  VGA_l074_g12468 : AOI22D0BWP7T port map(A1 => VGA_l074_n_166, A2 => y_pos_e4(4), B1 => VGA_l074_n_159, B2 => VGA_l074_n_11, ZN => VGA_l074_n_179);
  VGA_l074_g12469 : ND2D0BWP7T port map(A1 => VGA_l074_n_168, A2 => VGA_l074_n_171, ZN => VGA_l074_n_177);
  VGA_l074_g12470 : ND2D0BWP7T port map(A1 => VGA_l074_n_164, A2 => VGA_l074_n_140, ZN => VGA_l074_n_176);
  VGA_l074_g12471 : CKND1BWP7T port map(I => VGA_l074_n_174, ZN => VGA_l074_n_175);
  VGA_l074_g12472 : OAI211D0BWP7T port map(A1 => VGA_l074_n_96, A2 => VGA_l074_n_129, B => VGA_l074_n_153, C => VGA_l074_n_105, ZN => VGA_l074_n_173);
  VGA_l074_g12473 : ND3D0BWP7T port map(A1 => VGA_l074_n_154, A2 => VGA_l074_n_158, A3 => VGA_l074_n_115, ZN => VGA_l074_n_172);
  VGA_l074_g12474 : ND3D0BWP7T port map(A1 => VGA_l074_n_159, A2 => VGA_l074_n_102, A3 => VGA_l074_n_37, ZN => VGA_l074_n_174);
  VGA_l074_g12475 : CKND1BWP7T port map(I => VGA_l074_n_168, ZN => VGA_l074_n_169);
  VGA_l074_g12476 : ND2D0BWP7T port map(A1 => VGA_l074_n_156, A2 => VGA_l074_n_114, ZN => VGA_l074_n_171);
  VGA_l074_g12477 : AN2D1BWP7T port map(A1 => VGA_l074_n_154, A2 => VGA_l074_n_113, Z => VGA_l074_n_170);
  VGA_l074_g12478 : ND2D0BWP7T port map(A1 => VGA_l074_n_160, A2 => VGA_l074_n_113, ZN => VGA_l074_n_168);
  VGA_l074_g12479 : ND2D0BWP7T port map(A1 => VGA_l074_n_155, A2 => VGA_l074_n_114, ZN => VGA_l074_n_167);
  VGA_l074_g12480 : AOI221D0BWP7T port map(A1 => VGA_l074_n_125, A2 => VGA_l074_n_95, B1 => VGA_l074_n_45, B2 => VGA_l074_n_81, C => VGA_l074_n_152, ZN => VGA_l074_n_163);
  VGA_l074_g12481 : AN4D1BWP7T port map(A1 => VGA_l074_n_141, A2 => VGA_l074_n_103, A3 => VGA_l074_n_89, A4 => VGA_l074_n_0, Z => VGA_l074_n_162);
  VGA_l074_g12482 : NR3D0BWP7T port map(A1 => VGA_l074_n_149, A2 => VGA_l074_n_44, A3 => VGA_y(4), ZN => VGA_l074_n_166);
  VGA_l074_g12483 : IND3D0BWP7T port map(A1 => VGA_l074_n_127, B1 => VGA_l074_n_2, B2 => VGA_l074_n_158, ZN => VGA_l074_n_165);
  VGA_l074_g12484 : AN2D1BWP7T port map(A1 => VGA_l074_n_158, A2 => VGA_l074_n_116, Z => VGA_l074_n_164);
  VGA_l074_g12485 : IINR4D0BWP7T port map(A1 => VGA_l074_n_122, A2 => VGA_l074_n_69, B1 => VGA_l074_n_133, B2 => VGA_l074_n_77, ZN => VGA_l074_n_157);
  VGA_l074_g12486 : IND2D0BWP7T port map(A1 => VGA_l074_n_151, B1 => VGA_l074_n_150, ZN => VGA_l074_n_161);
  VGA_l074_g12487 : NR3D0BWP7T port map(A1 => VGA_l074_n_148, A2 => VGA_l074_n_87, A3 => VGA_l074_n_40, ZN => VGA_l074_n_160);
  VGA_l074_g12488 : INR2D0BWP7T port map(A1 => VGA_l074_n_44, B1 => VGA_l074_n_149, ZN => VGA_l074_n_159);
  VGA_l074_g12489 : AOI211D0BWP7T port map(A1 => VGA_l074_n_44, A2 => VGA_l074_n_34, B => VGA_l074_n_149, C => VGA_l074_n_98, ZN => VGA_l074_n_158);
  VGA_l074_g12490 : AOI22D0BWP7T port map(A1 => VGA_l074_n_146, A2 => VGA_l074_n_126, B1 => VGA_l074_n_45, B2 => VGA_l074_n_26, ZN => VGA_l074_n_153);
  VGA_l074_g12491 : OAI22D0BWP7T port map(A1 => VGA_l074_n_146, A2 => VGA_l074_n_130, B1 => VGA_l074_n_97, B2 => VGA_x(5), ZN => VGA_l074_n_152);
  VGA_l074_g12492 : INR3D0BWP7T port map(A1 => VGA_l074_n_148, B1 => VGA_l074_n_40, B2 => VGA_l074_n_87, ZN => VGA_l074_n_156);
  VGA_l074_g12493 : AN3D0BWP7T port map(A1 => VGA_l074_n_147, A2 => VGA_l074_n_87, A3 => VGA_l074_n_39, Z => VGA_l074_n_155);
  VGA_l074_g12494 : INR3D0BWP7T port map(A1 => VGA_l074_n_87, B1 => VGA_l074_n_40, B2 => VGA_l074_n_147, ZN => VGA_l074_n_154);
  VGA_l074_g12495 : AN2D1BWP7T port map(A1 => VGA_l074_n_144, A2 => VGA_l074_n_114, Z => VGA_l074_n_151);
  VGA_l074_g12496 : ND2D0BWP7T port map(A1 => VGA_l074_n_143, A2 => VGA_l074_n_113, ZN => VGA_l074_n_150);
  VGA_l074_g12497 : IND4D0BWP7T port map(A1 => VGA_l074_n_108, B1 => VGA_l074_n_109, B2 => VGA_l074_n_106, B3 => VGA_l074_n_107, ZN => VGA_l074_n_149);
  VGA_l074_g12498 : AN3D0BWP7T port map(A1 => VGA_l074_n_128, A2 => VGA_l074_n_70, A3 => VGA_l074_n_76, Z => VGA_l074_n_145);
  VGA_l074_g12499 : OAI221D0BWP7T port map(A1 => VGA_l074_n_101, A2 => y_pos_e4(1), B1 => VGA_l074_n_4, B2 => VGA_l074_n_82, C => VGA_l074_n_100, ZN => VGA_l074_n_148);
  VGA_l074_g12500 : OAI211D0BWP7T port map(A1 => y_pos_e4(1), A2 => VGA_l074_n_41, B => VGA_l074_n_121, C => VGA_l074_n_101, ZN => VGA_l074_n_147);
  VGA_l074_g12501 : MAOI222D0BWP7T port map(A => VGA_x(2), B => x_pos_e4(2), C => VGA_l074_n_83, ZN => VGA_l074_n_146);
  VGA_l074_g12502 : AN3D0BWP7T port map(A1 => VGA_l074_n_124, A2 => VGA_l074_n_94, A3 => VGA_l074_n_92, Z => VGA_l074_n_142);
  VGA_l074_g12503 : INR3D0BWP7T port map(A1 => VGA_l074_n_128, B1 => VGA_l074_n_72, B2 => VGA_l074_n_77, ZN => VGA_l074_n_141);
  VGA_l074_g12504 : AOI211D0BWP7T port map(A1 => VGA_l074_n_101, A2 => VGA_l074_n_100, B => VGA_l074_n_39, C => VGA_l074_n_43, ZN => VGA_l074_n_144);
  VGA_l074_g12505 : AN4D1BWP7T port map(A1 => VGA_l074_n_101, A2 => VGA_l074_n_100, A3 => VGA_l074_n_42, A4 => VGA_l074_n_40, Z => VGA_l074_n_143);
  VGA_l074_g12506 : INR2D0BWP7T port map(A1 => VGA_l074_n_122, B1 => VGA_l074_n_72, ZN => VGA_l074_n_139);
  VGA_l074_g12507 : AN2D1BWP7T port map(A1 => VGA_l074_n_112, A2 => VGA_l074_n_52, Z => VGA_l074_n_138);
  VGA_l074_g12508 : ND2D0BWP7T port map(A1 => VGA_l074_n_123, A2 => VGA_l074_n_131, ZN => VGA_l074_n_137);
  VGA_l074_g12509 : INR2D0BWP7T port map(A1 => VGA_l074_n_104, B1 => VGA_l074_n_1, ZN => VGA_l074_n_140);
  VGA_l074_g12510 : OA221D0BWP7T port map(A1 => VGA_l074_n_67, A2 => VGA_draw_count8(1), B1 => VGA_l074_n_24, B2 => VGA_l074_n_54, C => VGA_l074_n_74, Z => VGA_l074_n_135);
  VGA_l074_g12511 : OAI211D0BWP7T port map(A1 => VGA_draw_count8(1), A2 => VGA_l074_n_58, B => VGA_l074_n_84, C => VGA_l074_n_74, ZN => VGA_l074_n_134);
  VGA_l074_g12512 : OAI211D0BWP7T port map(A1 => VGA_l074_n_13, A2 => VGA_l074_n_54, B => VGA_l074_n_85, C => VGA_l074_n_75, ZN => VGA_l074_n_133);
  VGA_l074_g12513 : OA21D0BWP7T port map(A1 => VGA_l074_n_14, A2 => VGA_l074_n_3, B => VGA_l074_n_124, Z => VGA_l074_n_132);
  VGA_l074_g12514 : ND2D0BWP7T port map(A1 => VGA_l074_n_110, A2 => VGA_l074_n_105, ZN => VGA_l074_n_136);
  VGA_l074_g12515 : CKND1BWP7T port map(I => VGA_l074_n_129, ZN => VGA_l074_n_130);
  VGA_l074_g12516 : CKND1BWP7T port map(I => VGA_l074_n_125, ZN => VGA_l074_n_126);
  VGA_l074_g12517 : IND2D0BWP7T port map(A1 => VGA_l074_n_100, B1 => y_pos_e4(1), ZN => VGA_l074_n_121);
  VGA_l074_g12518 : MOAI22D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l074_n_10, B1 => VGA_l074_n_49, B2 => VGA_l074_n_32, ZN => VGA_l074_n_120);
  VGA_l074_g12519 : AOI21D0BWP7T port map(A1 => VGA_l074_n_59, A2 => VGA_l074_n_27, B => VGA_l074_n_93, ZN => VGA_l074_n_119);
  VGA_l074_g12520 : AOI211D0BWP7T port map(A1 => VGA_l074_n_55, A2 => VGA_l074_n_24, B => VGA_l074_n_93, C => VGA_l074_n_78, ZN => VGA_l074_n_118);
  VGA_l074_g12521 : OAI221D0BWP7T port map(A1 => VGA_l074_n_62, A2 => VGA_l074_n_0, B1 => VGA_l074_n_29, B2 => VGA_l074_n_64, C => VGA_l074_n_92, ZN => VGA_l074_n_117);
  VGA_l074_g12522 : OA21D0BWP7T port map(A1 => VGA_l074_n_62, A2 => VGA_l074_n_64, B => VGA_l074_n_92, Z => VGA_l074_n_131);
  VGA_l074_g12523 : AOI22D0BWP7T port map(A1 => VGA_l074_n_66, A2 => VGA_l074_n_31, B1 => VGA_l074_n_47, B2 => VGA_x(2), ZN => VGA_l074_n_129);
  VGA_l074_g12524 : NR3D0BWP7T port map(A1 => VGA_l074_n_80, A2 => VGA_l074_n_73, A3 => VGA_l074_n_61, ZN => VGA_l074_n_128);
  VGA_l074_g12525 : IND2D0BWP7T port map(A1 => VGA_l074_n_37, B1 => VGA_l074_n_102, ZN => VGA_l074_n_127);
  VGA_l074_g12526 : OAI22D0BWP7T port map(A1 => VGA_l074_n_66, A2 => VGA_l074_n_31, B1 => VGA_l074_n_47, B2 => VGA_x(2), ZN => VGA_l074_n_125);
  VGA_l074_g12527 : AN3D0BWP7T port map(A1 => VGA_l074_n_68, A2 => VGA_l074_n_75, A3 => VGA_l074_n_69, Z => VGA_l074_n_124);
  VGA_l074_g12528 : AN2D1BWP7T port map(A1 => VGA_l074_n_88, A2 => VGA_l074_n_68, Z => VGA_l074_n_123);
  VGA_l074_g12529 : AN2D1BWP7T port map(A1 => VGA_l074_n_89, A2 => VGA_l074_n_58, Z => VGA_l074_n_122);
  VGA_l074_g12530 : AOI221D0BWP7T port map(A1 => VGA_l074_n_61, A2 => VGA_draw_count8(0), B1 => VGA_l074_n_56, B2 => VGA_l074_n_25, C => VGA_l074_n_80, ZN => VGA_l074_n_112);
  VGA_l074_g12531 : AO222D0BWP7T port map(A1 => VGA_l074_n_61, A2 => VGA_l074_n_24, B1 => VGA_l074_n_55, B2 => VGA_l074_n_13, C1 => VGA_l074_n_53, C2 => VGA_l074_n_27, Z => VGA_l074_n_111);
  VGA_l074_g12532 : OAI22D0BWP7T port map(A1 => VGA_l074_n_45, A2 => VGA_l074_n_26, B1 => VGA_l074_n_46, B2 => VGA_l074_n_16, ZN => VGA_l074_n_110);
  VGA_l074_g12533 : MAOI22D0BWP7T port map(A1 => VGA_l074_n_50, A2 => VGA_l074_n_35, B1 => VGA_l074_n_50, B2 => VGA_l074_n_35, ZN => VGA_l074_n_109);
  VGA_l074_g12534 : OAI22D0BWP7T port map(A1 => VGA_l074_n_65, A2 => VGA_l074_n_15, B1 => VGA_l074_n_36, B2 => VGA_y(9), ZN => VGA_l074_n_108);
  VGA_l074_g12535 : AOI22D0BWP7T port map(A1 => VGA_l074_n_65, A2 => VGA_l074_n_15, B1 => VGA_l074_n_36, B2 => VGA_y(9), ZN => VGA_l074_n_107);
  VGA_l074_g12536 : MAOI22D0BWP7T port map(A1 => VGA_l074_n_48, A2 => VGA_l074_n_28, B1 => VGA_l074_n_48, B2 => VGA_l074_n_28, ZN => VGA_l074_n_106);
  VGA_l074_g12538 : MAOI22D0BWP7T port map(A1 => VGA_l074_n_38, A2 => VGA_l074_n_19, B1 => VGA_l074_n_38, B2 => VGA_l074_n_19, ZN => VGA_l074_n_116);
  VGA_l074_g12540 : MOAI22D0BWP7T port map(A1 => VGA_l074_n_38, A2 => VGA_l074_n_22, B1 => VGA_l074_n_38, B2 => VGA_l074_n_22, ZN => VGA_l074_n_115);
  VGA_l074_g12541 : MAOI22D0BWP7T port map(A1 => VGA_l074_n_37, A2 => VGA_l074_n_33, B1 => VGA_l074_n_37, B2 => VGA_l074_n_33, ZN => VGA_l074_n_114);
  VGA_l074_g12542 : MOAI22D0BWP7T port map(A1 => VGA_l074_n_37, A2 => VGA_l074_n_23, B1 => VGA_l074_n_37, B2 => VGA_l074_n_23, ZN => VGA_l074_n_113);
  VGA_l074_g12543 : AOI21D0BWP7T port map(A1 => VGA_l074_n_56, A2 => VGA_l074_n_24, B => VGA_l074_n_63, ZN => VGA_l074_n_99);
  VGA_l074_g12544 : NR2D0BWP7T port map(A1 => VGA_l074_n_44, A2 => VGA_l074_n_34, ZN => VGA_l074_n_98);
  VGA_l074_g12545 : IND2D0BWP7T port map(A1 => VGA_l074_n_46, B1 => x_pos_e4(5), ZN => VGA_l074_n_97);
  VGA_l074_g12546 : ND2D0BWP7T port map(A1 => VGA_l074_n_46, A2 => VGA_l074_n_16, ZN => VGA_l074_n_105);
  VGA_l074_g12547 : NR2D0BWP7T port map(A1 => VGA_l074_n_66, A2 => VGA_l074_n_31, ZN => VGA_l074_n_96);
  VGA_l074_g12548 : NR2D0BWP7T port map(A1 => VGA_l074_n_71, A2 => VGA_l074_n_41, ZN => VGA_l074_n_104);
  VGA_l074_g12550 : NR2D0BWP7T port map(A1 => VGA_l074_n_79, A2 => VGA_l074_n_78, ZN => VGA_l074_n_103);
  VGA_l074_g12551 : NR2D0BWP7T port map(A1 => VGA_l074_n_71, A2 => VGA_l074_n_82, ZN => VGA_l074_n_102);
  VGA_l074_g12552 : ND2D0BWP7T port map(A1 => VGA_l074_n_82, A2 => VGA_y(1), ZN => VGA_l074_n_101);
  VGA_l074_g12553 : IND2D0BWP7T port map(A1 => VGA_y(1), B1 => VGA_l074_n_41, ZN => VGA_l074_n_100);
  VGA_l074_g12554 : CKND1BWP7T port map(I => VGA_l074_n_90, ZN => VGA_l074_n_91);
  VGA_l074_g12555 : AOI21D0BWP7T port map(A1 => VGA_l074_n_59, A2 => VGA_l074_n_25, B => VGA_l074_n_73, ZN => VGA_l074_n_86);
  VGA_l074_g12556 : OAI21D0BWP7T port map(A1 => VGA_l074_n_56, A2 => VGA_l074_n_53, B => VGA_l074_n_24, ZN => VGA_l074_n_85);
  VGA_l074_g12557 : AO21D0BWP7T port map(A1 => VGA_l074_n_60, A2 => VGA_l074_n_54, B => VGA_l074_n_62, Z => VGA_l074_n_84);
  VGA_l074_g12558 : IAO21D0BWP7T port map(A1 => VGA_l074_n_60, A2 => VGA_l074_n_13, B => VGA_l074_n_55, ZN => VGA_l074_n_94);
  VGA_l074_g12559 : OAI21D0BWP7T port map(A1 => VGA_l074_n_52, A2 => VGA_draw_count8(1), B => VGA_l074_n_70, ZN => VGA_l074_n_93);
  VGA_l074_g12560 : AOI22D0BWP7T port map(A1 => VGA_l074_n_51, A2 => VGA_x(0), B1 => VGA_x(1), B2 => VGA_l074_n_6, ZN => VGA_l074_n_83);
  VGA_l074_g12561 : OA22D0BWP7T port map(A1 => VGA_l074_n_64, A2 => VGA_l074_n_12, B1 => VGA_l074_n_25, B2 => VGA_l074_n_0, Z => VGA_l074_n_92);
  VGA_l074_g12562 : OAI21D0BWP7T port map(A1 => VGA_l074_n_57, A2 => VGA_l074_n_13, B => VGA_l074_n_69, ZN => VGA_l074_n_90);
  VGA_l074_g12563 : AOI22D0BWP7T port map(A1 => VGA_l074_n_56, A2 => VGA_l074_n_13, B1 => VGA_l074_n_59, B2 => VGA_l074_n_24, ZN => VGA_l074_n_89);
  VGA_l074_g12564 : IAO21D0BWP7T port map(A1 => VGA_l074_n_0, A2 => VGA_l074_n_24, B => VGA_l074_n_79, ZN => VGA_l074_n_88);
  VGA_l074_g12565 : MOAI22D0BWP7T port map(A1 => VGA_l074_n_43, A2 => VGA_y(0), B1 => VGA_l074_n_43, B2 => VGA_y(0), ZN => VGA_l074_n_87);
  VGA_l074_g12568 : INVD0BWP7T port map(I => VGA_l074_n_41, ZN => VGA_l074_n_82);
  VGA_l074_g12569 : CKND1BWP7T port map(I => VGA_l074_n_26, ZN => VGA_l074_n_81);
  VGA_l074_g12570 : NR2D0BWP7T port map(A1 => VGA_l074_n_54, A2 => VGA_draw_count8(1), ZN => VGA_l074_n_80);
  VGA_l074_g12571 : INR2D0BWP7T port map(A1 => VGA_l074_n_63, B1 => VGA_l074_n_25, ZN => VGA_l074_n_79);
  VGA_l074_g12572 : NR2D0BWP7T port map(A1 => VGA_l074_n_0, A2 => VGA_draw_count8(1), ZN => VGA_l074_n_78);
  VGA_l074_g12573 : NR2D0BWP7T port map(A1 => VGA_l074_n_57, A2 => VGA_l074_n_29, ZN => VGA_l074_n_77);
  VGA_l074_g12574 : ND2D0BWP7T port map(A1 => VGA_l074_n_55, A2 => VGA_draw_count8(1), ZN => VGA_l074_n_76);
  VGA_l074_g12575 : ND2D0BWP7T port map(A1 => VGA_l074_n_53, A2 => VGA_l074_n_13, ZN => VGA_l074_n_75);
  VGA_l074_g12576 : ND2D0BWP7T port map(A1 => VGA_l074_n_53, A2 => VGA_draw_count8(1), ZN => VGA_l074_n_74);
  VGA_l074_g12577 : NR2D0BWP7T port map(A1 => VGA_l074_n_56, A2 => VGA_l074_n_59, ZN => VGA_l074_n_67);
  VGA_l074_g12578 : AN2D1BWP7T port map(A1 => VGA_l074_n_63, A2 => VGA_l074_n_27, Z => VGA_l074_n_73);
  VGA_l074_g12579 : NR2D0BWP7T port map(A1 => VGA_l074_n_52, A2 => VGA_l074_n_13, ZN => VGA_l074_n_72);
  VGA_l074_g12580 : ND2D0BWP7T port map(A1 => VGA_l074_n_40, A2 => VGA_l074_n_43, ZN => VGA_l074_n_71);
  VGA_l074_g12581 : IND2D0BWP7T port map(A1 => VGA_l074_n_62, B1 => VGA_l074_n_56, ZN => VGA_l074_n_70);
  VGA_l074_g12582 : ND2D0BWP7T port map(A1 => VGA_l074_n_63, A2 => VGA_l074_n_13, ZN => VGA_l074_n_69);
  VGA_l074_g12583 : IND2D0BWP7T port map(A1 => VGA_l074_n_62, B1 => VGA_l074_n_63, ZN => VGA_l074_n_68);
  VGA_l074_g12584 : INVD0BWP7T port map(I => VGA_l074_n_61, ZN => VGA_l074_n_60);
  VGA_l074_g12585 : INVD0BWP7T port map(I => VGA_l074_n_59, ZN => VGA_l074_n_58);
  VGA_l074_g12586 : INVD1BWP7T port map(I => VGA_l074_n_57, ZN => VGA_l074_n_56);
  VGA_l074_g12587 : INVD0BWP7T port map(I => VGA_l074_n_55, ZN => VGA_l074_n_54);
  VGA_l074_g12588 : INVD0BWP7T port map(I => VGA_l074_n_53, ZN => VGA_l074_n_52);
  VGA_l074_g12589 : IAO21D0BWP7T port map(A1 => VGA_x(1), A2 => VGA_l074_n_6, B => x_pos_e4(0), ZN => VGA_l074_n_51);
  VGA_l074_g12590 : OAI21D0BWP7T port map(A1 => VGA_l074_n_7, A2 => x_pos_e4(4), B => VGA_l074_n_26, ZN => VGA_l074_n_66);
  VGA_l074_g12591 : AOI21D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l074_n_5, B => VGA_l074_n_28, ZN => VGA_l074_n_65);
  VGA_l074_g12592 : IND2D0BWP7T port map(A1 => VGA_l074_n_30, B1 => VGA_draw_count8(4), ZN => VGA_l074_n_64);
  VGA_l074_g12593 : INR2D0BWP7T port map(A1 => VGA_draw_count8(4), B1 => VGA_l074_n_17, ZN => VGA_l074_n_63);
  VGA_l074_g12594 : INR2D0BWP7T port map(A1 => VGA_l074_n_29, B1 => VGA_l074_n_27, ZN => VGA_l074_n_62);
  VGA_l074_g12596 : NR2D0BWP7T port map(A1 => VGA_l074_n_14, A2 => VGA_draw_count8(4), ZN => VGA_l074_n_61);
  VGA_l074_g12597 : NR2D0BWP7T port map(A1 => VGA_l074_n_30, A2 => VGA_draw_count8(4), ZN => VGA_l074_n_59);
  VGA_l074_g12598 : IND2D0BWP7T port map(A1 => VGA_l074_n_14, B1 => VGA_draw_count8(4), ZN => VGA_l074_n_57);
  VGA_l074_g12599 : NR2D0BWP7T port map(A1 => VGA_l074_n_17, A2 => VGA_draw_count8(4), ZN => VGA_l074_n_55);
  VGA_l074_g12600 : NR2D0BWP7T port map(A1 => VGA_l074_n_18, A2 => VGA_draw_count8(4), ZN => VGA_l074_n_53);
  VGA_l074_g12601 : CKND1BWP7T port map(I => VGA_l074_n_43, ZN => VGA_l074_n_42);
  VGA_l074_g12602 : CKND1BWP7T port map(I => VGA_l074_n_40, ZN => VGA_l074_n_39);
  VGA_l074_g12603 : MOAI22D0BWP7T port map(A1 => VGA_y(8), A2 => y_pos_e4(8), B1 => VGA_y(8), B2 => y_pos_e4(8), ZN => VGA_l074_n_50);
  VGA_l074_g12604 : MOAI22D0BWP7T port map(A1 => VGA_x(7), A2 => x_pos_e4(7), B1 => VGA_x(7), B2 => x_pos_e4(7), ZN => VGA_l074_n_49);
  VGA_l074_g12605 : MOAI22D0BWP7T port map(A1 => VGA_y(7), A2 => y_pos_e4(7), B1 => VGA_y(7), B2 => y_pos_e4(7), ZN => VGA_l074_n_48);
  VGA_l074_g12606 : MAOI22D0BWP7T port map(A1 => VGA_x(3), A2 => x_pos_e4(3), B1 => VGA_x(3), B2 => x_pos_e4(3), ZN => VGA_l074_n_47);
  VGA_l074_g12607 : MOAI22D0BWP7T port map(A1 => VGA_x(6), A2 => x_pos_e4(6), B1 => VGA_x(6), B2 => x_pos_e4(6), ZN => VGA_l074_n_46);
  VGA_l074_g12608 : MOAI22D0BWP7T port map(A1 => VGA_x(5), A2 => x_pos_e4(5), B1 => VGA_x(5), B2 => x_pos_e4(5), ZN => VGA_l074_n_45);
  VGA_l074_g12609 : MAOI22D0BWP7T port map(A1 => VGA_y(5), A2 => y_pos_e4(5), B1 => VGA_y(5), B2 => y_pos_e4(5), ZN => VGA_l074_n_44);
  VGA_l074_g12610 : MOAI22D0BWP7T port map(A1 => VGA_y(1), A2 => y_pos_e4(1), B1 => VGA_y(1), B2 => y_pos_e4(1), ZN => VGA_l074_n_43);
  VGA_l074_g12611 : MOAI22D0BWP7T port map(A1 => VGA_y(2), A2 => y_pos_e4(2), B1 => VGA_y(2), B2 => y_pos_e4(2), ZN => VGA_l074_n_41);
  VGA_l074_g12612 : MOAI22D0BWP7T port map(A1 => VGA_y(0), A2 => y_pos_e4(0), B1 => VGA_y(0), B2 => y_pos_e4(0), ZN => VGA_l074_n_40);
  VGA_l074_g12613 : MAOI22D0BWP7T port map(A1 => VGA_y(4), A2 => y_pos_e4(4), B1 => VGA_y(4), B2 => y_pos_e4(4), ZN => VGA_l074_n_38);
  VGA_l074_g12614 : MOAI22D0BWP7T port map(A1 => VGA_y(3), A2 => y_pos_e4(3), B1 => VGA_y(3), B2 => y_pos_e4(3), ZN => VGA_l074_n_37);
  VGA_l074_g12615 : INVD1BWP7T port map(I => VGA_l074_n_25, ZN => VGA_l074_n_24);
  VGA_l074_g12616 : IND2D0BWP7T port map(A1 => VGA_y(8), B1 => y_pos_e4(8), ZN => VGA_l074_n_36);
  VGA_l074_g12617 : INR2D0BWP7T port map(A1 => y_pos_e4(7), B1 => VGA_y(7), ZN => VGA_l074_n_35);
  VGA_l074_g12618 : IND2D0BWP7T port map(A1 => y_pos_e4(4), B1 => VGA_y(4), ZN => VGA_l074_n_34);
  VGA_l074_g12619 : IND2D0BWP7T port map(A1 => y_pos_e4(2), B1 => VGA_y(2), ZN => VGA_l074_n_33);
  VGA_l074_g12620 : IND2D0BWP7T port map(A1 => x_pos_e4(6), B1 => VGA_x(6), ZN => VGA_l074_n_32);
  VGA_l074_g12621 : IND2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_e4(3), ZN => VGA_l074_n_31);
  VGA_l074_g12622 : ND2D0BWP7T port map(A1 => VGA_draw_count8(2), A2 => VGA_draw_count8(3), ZN => VGA_l074_n_30);
  VGA_l074_g12623 : ND2D0BWP7T port map(A1 => VGA_l074_n_3, A2 => VGA_draw_count8(0), ZN => VGA_l074_n_29);
  VGA_l074_g12624 : NR2D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l074_n_5, ZN => VGA_l074_n_28);
  VGA_l074_g12625 : NR2D0BWP7T port map(A1 => VGA_l074_n_3, A2 => VGA_draw_count8(0), ZN => VGA_l074_n_27);
  VGA_l074_g12626 : ND2D0BWP7T port map(A1 => VGA_l074_n_7, A2 => x_pos_e4(4), ZN => VGA_l074_n_26);
  VGA_l074_g12627 : ND2D0BWP7T port map(A1 => VGA_draw_count8(1), A2 => VGA_draw_count8(0), ZN => VGA_l074_n_25);
  VGA_l074_g12629 : CKND1BWP7T port map(I => VGA_l074_n_13, ZN => VGA_l074_n_12);
  VGA_l074_g12630 : IND2D0BWP7T port map(A1 => VGA_y(4), B1 => y_pos_e4(4), ZN => VGA_l074_n_11);
  VGA_l074_g12631 : ND2D0BWP7T port map(A1 => VGA_l074_n_8, A2 => y_pos_e4(2), ZN => VGA_l074_n_23);
  VGA_l074_g12632 : NR2D0BWP7T port map(A1 => VGA_l074_n_9, A2 => y_pos_e4(3), ZN => VGA_l074_n_22);
  VGA_l074_g12633 : INR2D0BWP7T port map(A1 => x_pos_e4(7), B1 => VGA_x(7), ZN => VGA_l074_n_21);
  VGA_l074_g12634 : ND2D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l074_n_10, ZN => VGA_l074_n_20);
  VGA_l074_g12635 : INR2D0BWP7T port map(A1 => y_pos_e4(3), B1 => VGA_y(3), ZN => VGA_l074_n_19);
  VGA_l074_g12636 : IND2D0BWP7T port map(A1 => VGA_draw_count8(2), B1 => VGA_draw_count8(3), ZN => VGA_l074_n_18);
  VGA_l074_g12637 : IND2D0BWP7T port map(A1 => VGA_draw_count8(3), B1 => VGA_draw_count8(2), ZN => VGA_l074_n_17);
  VGA_l074_g12638 : INR2D0BWP7T port map(A1 => VGA_x(5), B1 => x_pos_e4(5), ZN => VGA_l074_n_16);
  VGA_l074_g12639 : IND2D0BWP7T port map(A1 => y_pos_e4(5), B1 => VGA_y(5), ZN => VGA_l074_n_15);
  VGA_l074_g12640 : OR2D0BWP7T port map(A1 => VGA_draw_count8(2), A2 => VGA_draw_count8(3), Z => VGA_l074_n_14);
  VGA_l074_g12641 : NR2D0BWP7T port map(A1 => VGA_draw_count8(1), A2 => VGA_draw_count8(0), ZN => VGA_l074_n_13);
  VGA_l074_g12642 : CKND1BWP7T port map(I => x_pos_e4(8), ZN => VGA_l074_n_10);
  VGA_l074_g12643 : CKND1BWP7T port map(I => VGA_y(3), ZN => VGA_l074_n_9);
  VGA_l074_g12644 : CKND1BWP7T port map(I => VGA_y(2), ZN => VGA_l074_n_8);
  VGA_l074_g12645 : CKND1BWP7T port map(I => VGA_x(4), ZN => VGA_l074_n_7);
  VGA_l074_g12646 : CKND1BWP7T port map(I => x_pos_e4(1), ZN => VGA_l074_n_6);
  VGA_l074_g12647 : CKND1BWP7T port map(I => y_pos_e4(6), ZN => VGA_l074_n_5);
  VGA_l074_g12648 : CKND1BWP7T port map(I => y_pos_e4(1), ZN => VGA_l074_n_4);
  VGA_l074_g12649 : INVD0BWP7T port map(I => VGA_draw_count8(1), ZN => VGA_l074_n_3);
  VGA_l074_g2 : MUX2ND0BWP7T port map(I0 => VGA_y(3), I1 => VGA_l074_n_9, S => VGA_l074_n_38, ZN => VGA_l074_n_2);
  VGA_l074_g12650 : MUX2ND0BWP7T port map(I0 => VGA_l074_n_8, I1 => VGA_y(2), S => VGA_l074_n_37, ZN => VGA_l074_n_1);
  VGA_l074_g12651 : IND2D1BWP7T port map(A1 => VGA_l074_n_18, B1 => VGA_draw_count8(4), ZN => VGA_l074_n_0);
  VGA_l074_g12652 : INVD0BWP7T port map(I => VGA_l074_n_66, ZN => VGA_l074_n_95);
  VGA_l075_g12402 : OAI211D0BWP7T port map(A1 => VGA_l075_n_76, A2 => VGA_l075_n_195, B => VGA_l075_n_243, C => VGA_l075_n_223, ZN => VGA_r9);
  VGA_l075_g12403 : AOI211D0BWP7T port map(A1 => VGA_l075_n_206, A2 => VGA_l075_n_111, B => VGA_l075_n_242, C => VGA_l075_n_225, ZN => VGA_l075_n_243);
  VGA_l075_g12404 : OAI211D0BWP7T port map(A1 => VGA_l075_n_162, A2 => VGA_l075_n_216, B => VGA_l075_n_241, C => VGA_l075_n_238, ZN => VGA_l075_n_242);
  VGA_l075_g12405 : NR4D0BWP7T port map(A1 => VGA_l075_n_239, A2 => VGA_l075_n_227, A3 => VGA_l075_n_219, A4 => VGA_l075_n_220, ZN => VGA_l075_n_241);
  VGA_l075_g12406 : OAI211D0BWP7T port map(A1 => VGA_l075_n_91, A2 => VGA_l075_n_212, B => VGA_l075_n_237, C => VGA_l075_n_235, ZN => VGA_g9);
  VGA_l075_g12407 : NR4D0BWP7T port map(A1 => VGA_l075_n_233, A2 => VGA_l075_n_191, A3 => VGA_l075_n_151, A4 => VGA_l075_n_138, ZN => VGA_l075_n_239);
  VGA_l075_g12408 : NR4D0BWP7T port map(A1 => VGA_l075_n_226, A2 => VGA_l075_n_228, A3 => VGA_l075_n_221, A4 => VGA_l075_n_192, ZN => VGA_l075_n_238);
  VGA_l075_g12409 : AOI211D0BWP7T port map(A1 => VGA_l075_n_206, A2 => VGA_l075_n_117, B => VGA_l075_n_236, C => VGA_l075_n_218, ZN => VGA_l075_n_237);
  VGA_l075_g12410 : OAI211D0BWP7T port map(A1 => VGA_l075_n_99, A2 => VGA_l075_n_195, B => VGA_l075_n_230, C => VGA_l075_n_224, ZN => VGA_l075_n_236);
  VGA_l075_g12411 : AOI211D0BWP7T port map(A1 => VGA_l075_n_211, A2 => VGA_l075_n_137, B => VGA_l075_n_231, C => VGA_l075_n_213, ZN => VGA_l075_n_235);
  VGA_l075_g12412 : OAI32D0BWP7T port map(A1 => VGA_l075_n_24, A2 => VGA_l075_n_60, A3 => VGA_l075_n_216, B1 => VGA_l075_n_94, B2 => VGA_l075_n_215, ZN => VGA_b9);
  VGA_l075_g12413 : ND4D0BWP7T port map(A1 => VGA_l075_n_210, A2 => VGA_l075_n_189, A3 => VGA_l075_n_176, A4 => VGA_l075_n_165, ZN => VGA_l075_n_233);
  VGA_l075_g12414 : OAI211D0BWP7T port map(A1 => VGA_l075_n_191, A2 => VGA_l075_n_209, B => VGA_l075_n_204, C => VGA_l075_n_199, ZN => VGA_enable9);
  VGA_l075_g12415 : OAI22D0BWP7T port map(A1 => VGA_l075_n_217, A2 => VGA_l075_n_139, B1 => VGA_l075_n_207, B2 => VGA_l075_n_131, ZN => VGA_l075_n_231);
  VGA_l075_g12416 : AOI31D0BWP7T port map(A1 => VGA_l075_n_190, A2 => VGA_l075_n_182, A3 => VGA_l075_n_77, B => VGA_l075_n_229, ZN => VGA_l075_n_230);
  VGA_l075_g12417 : AOI21D0BWP7T port map(A1 => VGA_l075_n_103, A2 => VGA_l075_n_86, B => VGA_l075_n_216, ZN => VGA_l075_n_229);
  VGA_l075_g12418 : AOI31D0BWP7T port map(A1 => VGA_l075_n_145, A2 => VGA_l075_n_88, A3 => VGA_l075_n_75, B => VGA_l075_n_217, ZN => VGA_l075_n_228);
  VGA_l075_g12419 : AOI31D0BWP7T port map(A1 => VGA_l075_n_122, A2 => VGA_l075_n_118, A3 => VGA_l075_n_60, B => VGA_l075_n_214, ZN => VGA_l075_n_227);
  VGA_l075_g12420 : AOI31D0BWP7T port map(A1 => VGA_l075_n_142, A2 => VGA_l075_n_122, A3 => VGA_l075_n_88, B => VGA_l075_n_215, ZN => VGA_l075_n_226);
  VGA_l075_g12421 : AOI22D0BWP7T port map(A1 => VGA_l075_n_205, A2 => VGA_l075_n_195, B1 => VGA_l075_n_119, B2 => VGA_l075_n_89, ZN => VGA_l075_n_225);
  VGA_l075_g12422 : AO21D0BWP7T port map(A1 => VGA_l075_n_123, A2 => VGA_l075_n_91, B => VGA_l075_n_215, Z => VGA_l075_n_224);
  VGA_l075_g12423 : OA21D0BWP7T port map(A1 => VGA_l075_n_208, A2 => VGA_l075_n_157, B => VGA_l075_n_222, Z => VGA_l075_n_223);
  VGA_l075_g12424 : AO31D0BWP7T port map(A1 => VGA_l075_n_135, A2 => VGA_l075_n_68, A3 => VGA_l075_n_69, B => VGA_l075_n_204, Z => VGA_l075_n_222);
  VGA_l075_g12425 : AOI21D0BWP7T port map(A1 => VGA_l075_n_89, A2 => VGA_l075_n_52, B => VGA_l075_n_212, ZN => VGA_l075_n_221);
  VGA_l075_g12426 : AOI31D0BWP7T port map(A1 => VGA_l075_n_132, A2 => VGA_l075_n_76, A3 => VGA_l075_n_58, B => VGA_l075_n_207, ZN => VGA_l075_n_220);
  VGA_l075_g12427 : OA21D0BWP7T port map(A1 => VGA_l075_n_134, A2 => VGA_l075_n_90, B => VGA_l075_n_211, Z => VGA_l075_n_219);
  VGA_l075_g12428 : AOI21D0BWP7T port map(A1 => VGA_l075_n_88, A2 => VGA_l075_n_0, B => VGA_l075_n_204, ZN => VGA_l075_n_218);
  VGA_l075_g12429 : AOI32D0BWP7T port map(A1 => VGA_l075_n_190, A2 => VGA_l075_n_181, A3 => VGA_l075_n_38, B1 => VGA_l075_n_202, B2 => VGA_l075_n_154, ZN => VGA_l075_n_214);
  VGA_l075_g12430 : AOI21D0BWP7T port map(A1 => VGA_l075_n_103, A2 => VGA_l075_n_68, B => VGA_l075_n_208, ZN => VGA_l075_n_213);
  VGA_l075_g12431 : AOI22D0BWP7T port map(A1 => VGA_l075_n_203, A2 => VGA_l075_n_156, B1 => VGA_l075_n_202, B2 => VGA_l075_n_143, ZN => VGA_l075_n_217);
  VGA_l075_g12432 : AOI22D0BWP7T port map(A1 => VGA_l075_n_202, A2 => VGA_l075_n_160, B1 => VGA_l075_n_203, B2 => VGA_l075_n_144, ZN => VGA_l075_n_216);
  VGA_l075_g12433 : AOI32D0BWP7T port map(A1 => VGA_l075_n_198, A2 => VGA_l075_n_1, A3 => VGA_l075_n_104, B1 => VGA_l075_n_203, B2 => VGA_l075_n_155, ZN => VGA_l075_n_215);
  VGA_l075_g12434 : OAI31D0BWP7T port map(A1 => VGA_l075_n_2, A2 => VGA_l075_n_127, A3 => VGA_l075_n_179, B => VGA_l075_n_201, ZN => VGA_l075_n_210);
  VGA_l075_g12435 : NR4D0BWP7T port map(A1 => VGA_l075_n_200, A2 => VGA_l075_n_186, A3 => VGA_l075_n_182, A4 => VGA_l075_n_185, ZN => VGA_l075_n_209);
  VGA_l075_g12436 : MAOI22D0BWP7T port map(A1 => VGA_l075_n_196, A2 => VGA_l075_n_170, B1 => VGA_l075_n_191, B2 => VGA_l075_n_165, ZN => VGA_l075_n_212);
  VGA_l075_g12437 : OAI22D0BWP7T port map(A1 => VGA_l075_n_197, A2 => VGA_l075_n_171, B1 => VGA_l075_n_193, B2 => VGA_l075_n_150, ZN => VGA_l075_n_211);
  VGA_l075_g12438 : CKND1BWP7T port map(I => VGA_l075_n_206, ZN => VGA_l075_n_205);
  VGA_l075_g12439 : AOI22D0BWP7T port map(A1 => VGA_l075_n_196, A2 => VGA_l075_n_169, B1 => VGA_l075_n_194, B2 => VGA_l075_n_151, ZN => VGA_l075_n_208);
  VGA_l075_g12440 : MAOI22D0BWP7T port map(A1 => VGA_l075_n_196, A2 => VGA_l075_n_151, B1 => VGA_l075_n_193, B2 => VGA_l075_n_168, ZN => VGA_l075_n_207);
  VGA_l075_g12441 : OAI22D0BWP7T port map(A1 => VGA_l075_n_197, A2 => VGA_l075_n_167, B1 => VGA_l075_n_191, B2 => VGA_l075_n_176, ZN => VGA_l075_n_206);
  VGA_l075_g12442 : MAOI22D0BWP7T port map(A1 => VGA_l075_n_196, A2 => VGA_l075_n_140, B1 => VGA_l075_n_193, B2 => VGA_l075_n_167, ZN => VGA_l075_n_204);
  VGA_l075_g12443 : INR2D0BWP7T port map(A1 => VGA_l075_n_198, B1 => VGA_l075_n_114, ZN => VGA_l075_n_203);
  VGA_l075_g12444 : INR2D0BWP7T port map(A1 => VGA_l075_n_198, B1 => VGA_l075_n_113, ZN => VGA_l075_n_202);
  VGA_l075_g12445 : CKND1BWP7T port map(I => VGA_l075_n_200, ZN => VGA_l075_n_201);
  VGA_l075_g12446 : OAI21D0BWP7T port map(A1 => VGA_l075_n_177, A2 => VGA_l075_n_161, B => VGA_l075_n_194, ZN => VGA_l075_n_199);
  VGA_l075_g12447 : ND3D0BWP7T port map(A1 => VGA_l075_n_188, A2 => VGA_l075_n_176, A3 => VGA_l075_n_165, ZN => VGA_l075_n_200);
  VGA_l075_g12448 : INVD0BWP7T port map(I => VGA_l075_n_197, ZN => VGA_l075_n_196);
  VGA_l075_g12449 : INR2D0BWP7T port map(A1 => VGA_l075_n_185, B1 => VGA_l075_n_191, ZN => VGA_l075_n_198);
  VGA_l075_g12450 : ND2D0BWP7T port map(A1 => VGA_l075_n_190, A2 => VGA_l075_n_184, ZN => VGA_l075_n_197);
  VGA_l075_g12451 : CKND1BWP7T port map(I => VGA_l075_n_193, ZN => VGA_l075_n_194);
  VGA_l075_g12452 : AOI211D0BWP7T port map(A1 => VGA_l075_n_122, A2 => VGA_l075_n_74, B => VGA_l075_n_191, C => VGA_l075_n_183, ZN => VGA_l075_n_192);
  VGA_l075_g12453 : IND2D0BWP7T port map(A1 => VGA_l075_n_189, B1 => VGA_l075_n_190, ZN => VGA_l075_n_195);
  VGA_l075_g12454 : ND2D0BWP7T port map(A1 => VGA_l075_n_190, A2 => VGA_l075_n_164, ZN => VGA_l075_n_193);
  VGA_l075_g12455 : INVD1BWP7T port map(I => VGA_l075_n_191, ZN => VGA_l075_n_190);
  VGA_l075_g12456 : OAI221D0BWP7T port map(A1 => VGA_l075_n_49, A2 => VGA_l075_n_32, B1 => VGA_l075_n_20, B2 => VGA_l075_n_21, C => VGA_l075_n_187, ZN => VGA_l075_n_191);
  VGA_l075_g12457 : AOI22D0BWP7T port map(A1 => VGA_l075_n_184, A2 => VGA_l075_n_161, B1 => VGA_l075_n_170, B2 => VGA_l075_n_164, ZN => VGA_l075_n_188);
  VGA_l075_g12458 : AOI33D0BWP7T port map(A1 => VGA_l075_n_184, A2 => VGA_l075_n_143, A3 => VGA_l075_n_113, B1 => VGA_l075_n_164, B2 => VGA_l075_n_156, B3 => VGA_l075_n_114, ZN => VGA_l075_n_189);
  VGA_l075_g12459 : AOI211D0BWP7T port map(A1 => VGA_l075_n_173, A2 => VGA_l075_n_136, B => VGA_l075_n_178, C => VGA_l075_n_120, ZN => VGA_l075_n_187);
  VGA_l075_g12460 : OA21D0BWP7T port map(A1 => VGA_l075_n_180, A2 => VGA_l075_n_170, B => VGA_l075_n_184, Z => VGA_l075_n_186);
  VGA_l075_g12461 : NR2D0BWP7T port map(A1 => VGA_l075_n_179, A2 => VGA_l075_n_115, ZN => VGA_l075_n_185);
  VGA_l075_g12462 : NR2D0BWP7T port map(A1 => VGA_l075_n_179, A2 => VGA_l075_n_116, ZN => VGA_l075_n_184);
  VGA_l075_g12463 : CKND1BWP7T port map(I => VGA_l075_n_182, ZN => VGA_l075_n_183);
  VGA_l075_g12464 : AO32D0BWP7T port map(A1 => VGA_l075_n_166, A2 => VGA_l075_n_102, A3 => VGA_l075_n_37, B1 => VGA_l075_n_175, B2 => VGA_y(4), Z => VGA_l075_n_181);
  VGA_l075_g12465 : OAI22D0BWP7T port map(A1 => VGA_l075_n_172, A2 => VGA_l075_n_113, B1 => VGA_l075_n_174, B2 => VGA_l075_n_38, ZN => VGA_l075_n_182);
  VGA_l075_g12466 : IND2D0BWP7T port map(A1 => VGA_l075_n_177, B1 => VGA_l075_n_167, ZN => VGA_l075_n_180);
  VGA_l075_g12467 : MOAI22D0BWP7T port map(A1 => VGA_l075_n_163, A2 => VGA_l075_n_136, B1 => VGA_l075_n_21, B2 => VGA_l075_n_20, ZN => VGA_l075_n_178);
  VGA_l075_g12468 : AOI22D0BWP7T port map(A1 => VGA_l075_n_166, A2 => y_pos_e5(4), B1 => VGA_l075_n_159, B2 => VGA_l075_n_11, ZN => VGA_l075_n_179);
  VGA_l075_g12469 : ND2D0BWP7T port map(A1 => VGA_l075_n_168, A2 => VGA_l075_n_171, ZN => VGA_l075_n_177);
  VGA_l075_g12470 : ND2D0BWP7T port map(A1 => VGA_l075_n_164, A2 => VGA_l075_n_140, ZN => VGA_l075_n_176);
  VGA_l075_g12471 : CKND1BWP7T port map(I => VGA_l075_n_174, ZN => VGA_l075_n_175);
  VGA_l075_g12472 : OAI211D0BWP7T port map(A1 => VGA_l075_n_96, A2 => VGA_l075_n_129, B => VGA_l075_n_153, C => VGA_l075_n_105, ZN => VGA_l075_n_173);
  VGA_l075_g12473 : ND3D0BWP7T port map(A1 => VGA_l075_n_154, A2 => VGA_l075_n_158, A3 => VGA_l075_n_115, ZN => VGA_l075_n_172);
  VGA_l075_g12474 : ND3D0BWP7T port map(A1 => VGA_l075_n_159, A2 => VGA_l075_n_102, A3 => VGA_l075_n_37, ZN => VGA_l075_n_174);
  VGA_l075_g12475 : CKND1BWP7T port map(I => VGA_l075_n_168, ZN => VGA_l075_n_169);
  VGA_l075_g12476 : ND2D0BWP7T port map(A1 => VGA_l075_n_156, A2 => VGA_l075_n_114, ZN => VGA_l075_n_171);
  VGA_l075_g12477 : AN2D1BWP7T port map(A1 => VGA_l075_n_154, A2 => VGA_l075_n_113, Z => VGA_l075_n_170);
  VGA_l075_g12478 : ND2D0BWP7T port map(A1 => VGA_l075_n_160, A2 => VGA_l075_n_113, ZN => VGA_l075_n_168);
  VGA_l075_g12479 : ND2D0BWP7T port map(A1 => VGA_l075_n_155, A2 => VGA_l075_n_114, ZN => VGA_l075_n_167);
  VGA_l075_g12480 : AOI221D0BWP7T port map(A1 => VGA_l075_n_125, A2 => VGA_l075_n_95, B1 => VGA_l075_n_45, B2 => VGA_l075_n_81, C => VGA_l075_n_152, ZN => VGA_l075_n_163);
  VGA_l075_g12481 : AN4D1BWP7T port map(A1 => VGA_l075_n_141, A2 => VGA_l075_n_103, A3 => VGA_l075_n_89, A4 => VGA_l075_n_0, Z => VGA_l075_n_162);
  VGA_l075_g12482 : NR3D0BWP7T port map(A1 => VGA_l075_n_149, A2 => VGA_l075_n_44, A3 => VGA_y(4), ZN => VGA_l075_n_166);
  VGA_l075_g12483 : IND3D0BWP7T port map(A1 => VGA_l075_n_127, B1 => VGA_l075_n_2, B2 => VGA_l075_n_158, ZN => VGA_l075_n_165);
  VGA_l075_g12484 : AN2D1BWP7T port map(A1 => VGA_l075_n_158, A2 => VGA_l075_n_116, Z => VGA_l075_n_164);
  VGA_l075_g12485 : IINR4D0BWP7T port map(A1 => VGA_l075_n_122, A2 => VGA_l075_n_69, B1 => VGA_l075_n_133, B2 => VGA_l075_n_77, ZN => VGA_l075_n_157);
  VGA_l075_g12486 : IND2D0BWP7T port map(A1 => VGA_l075_n_151, B1 => VGA_l075_n_150, ZN => VGA_l075_n_161);
  VGA_l075_g12487 : NR3D0BWP7T port map(A1 => VGA_l075_n_148, A2 => VGA_l075_n_87, A3 => VGA_l075_n_40, ZN => VGA_l075_n_160);
  VGA_l075_g12488 : INR2D0BWP7T port map(A1 => VGA_l075_n_44, B1 => VGA_l075_n_149, ZN => VGA_l075_n_159);
  VGA_l075_g12489 : AOI211D0BWP7T port map(A1 => VGA_l075_n_44, A2 => VGA_l075_n_34, B => VGA_l075_n_149, C => VGA_l075_n_98, ZN => VGA_l075_n_158);
  VGA_l075_g12490 : AOI22D0BWP7T port map(A1 => VGA_l075_n_146, A2 => VGA_l075_n_126, B1 => VGA_l075_n_45, B2 => VGA_l075_n_26, ZN => VGA_l075_n_153);
  VGA_l075_g12491 : OAI22D0BWP7T port map(A1 => VGA_l075_n_146, A2 => VGA_l075_n_130, B1 => VGA_l075_n_97, B2 => VGA_x(5), ZN => VGA_l075_n_152);
  VGA_l075_g12492 : INR3D0BWP7T port map(A1 => VGA_l075_n_148, B1 => VGA_l075_n_40, B2 => VGA_l075_n_87, ZN => VGA_l075_n_156);
  VGA_l075_g12493 : AN3D0BWP7T port map(A1 => VGA_l075_n_147, A2 => VGA_l075_n_87, A3 => VGA_l075_n_39, Z => VGA_l075_n_155);
  VGA_l075_g12494 : INR3D0BWP7T port map(A1 => VGA_l075_n_87, B1 => VGA_l075_n_40, B2 => VGA_l075_n_147, ZN => VGA_l075_n_154);
  VGA_l075_g12495 : AN2D1BWP7T port map(A1 => VGA_l075_n_144, A2 => VGA_l075_n_114, Z => VGA_l075_n_151);
  VGA_l075_g12496 : ND2D0BWP7T port map(A1 => VGA_l075_n_143, A2 => VGA_l075_n_113, ZN => VGA_l075_n_150);
  VGA_l075_g12497 : IND4D0BWP7T port map(A1 => VGA_l075_n_108, B1 => VGA_l075_n_109, B2 => VGA_l075_n_106, B3 => VGA_l075_n_107, ZN => VGA_l075_n_149);
  VGA_l075_g12498 : AN3D0BWP7T port map(A1 => VGA_l075_n_128, A2 => VGA_l075_n_70, A3 => VGA_l075_n_76, Z => VGA_l075_n_145);
  VGA_l075_g12499 : OAI221D0BWP7T port map(A1 => VGA_l075_n_101, A2 => y_pos_e5(1), B1 => VGA_l075_n_4, B2 => VGA_l075_n_82, C => VGA_l075_n_100, ZN => VGA_l075_n_148);
  VGA_l075_g12500 : OAI211D0BWP7T port map(A1 => y_pos_e5(1), A2 => VGA_l075_n_41, B => VGA_l075_n_121, C => VGA_l075_n_101, ZN => VGA_l075_n_147);
  VGA_l075_g12501 : MAOI222D0BWP7T port map(A => VGA_x(2), B => x_pos_e5(2), C => VGA_l075_n_83, ZN => VGA_l075_n_146);
  VGA_l075_g12502 : AN3D0BWP7T port map(A1 => VGA_l075_n_124, A2 => VGA_l075_n_94, A3 => VGA_l075_n_92, Z => VGA_l075_n_142);
  VGA_l075_g12503 : INR3D0BWP7T port map(A1 => VGA_l075_n_128, B1 => VGA_l075_n_72, B2 => VGA_l075_n_77, ZN => VGA_l075_n_141);
  VGA_l075_g12504 : AOI211D0BWP7T port map(A1 => VGA_l075_n_101, A2 => VGA_l075_n_100, B => VGA_l075_n_39, C => VGA_l075_n_43, ZN => VGA_l075_n_144);
  VGA_l075_g12505 : AN4D1BWP7T port map(A1 => VGA_l075_n_101, A2 => VGA_l075_n_100, A3 => VGA_l075_n_42, A4 => VGA_l075_n_40, Z => VGA_l075_n_143);
  VGA_l075_g12506 : INR2D0BWP7T port map(A1 => VGA_l075_n_122, B1 => VGA_l075_n_72, ZN => VGA_l075_n_139);
  VGA_l075_g12507 : AN2D1BWP7T port map(A1 => VGA_l075_n_112, A2 => VGA_l075_n_52, Z => VGA_l075_n_138);
  VGA_l075_g12508 : ND2D0BWP7T port map(A1 => VGA_l075_n_123, A2 => VGA_l075_n_131, ZN => VGA_l075_n_137);
  VGA_l075_g12509 : INR2D0BWP7T port map(A1 => VGA_l075_n_104, B1 => VGA_l075_n_1, ZN => VGA_l075_n_140);
  VGA_l075_g12510 : OA221D0BWP7T port map(A1 => VGA_l075_n_67, A2 => VGA_draw_count9(1), B1 => VGA_l075_n_24, B2 => VGA_l075_n_54, C => VGA_l075_n_74, Z => VGA_l075_n_135);
  VGA_l075_g12511 : OAI211D0BWP7T port map(A1 => VGA_draw_count9(1), A2 => VGA_l075_n_58, B => VGA_l075_n_84, C => VGA_l075_n_74, ZN => VGA_l075_n_134);
  VGA_l075_g12512 : OAI211D0BWP7T port map(A1 => VGA_l075_n_13, A2 => VGA_l075_n_54, B => VGA_l075_n_85, C => VGA_l075_n_75, ZN => VGA_l075_n_133);
  VGA_l075_g12513 : OA21D0BWP7T port map(A1 => VGA_l075_n_14, A2 => VGA_l075_n_3, B => VGA_l075_n_124, Z => VGA_l075_n_132);
  VGA_l075_g12514 : ND2D0BWP7T port map(A1 => VGA_l075_n_110, A2 => VGA_l075_n_105, ZN => VGA_l075_n_136);
  VGA_l075_g12515 : CKND1BWP7T port map(I => VGA_l075_n_129, ZN => VGA_l075_n_130);
  VGA_l075_g12516 : CKND1BWP7T port map(I => VGA_l075_n_125, ZN => VGA_l075_n_126);
  VGA_l075_g12517 : IND2D0BWP7T port map(A1 => VGA_l075_n_100, B1 => y_pos_e5(1), ZN => VGA_l075_n_121);
  VGA_l075_g12518 : MOAI22D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l075_n_10, B1 => VGA_l075_n_49, B2 => VGA_l075_n_32, ZN => VGA_l075_n_120);
  VGA_l075_g12519 : AOI21D0BWP7T port map(A1 => VGA_l075_n_59, A2 => VGA_l075_n_27, B => VGA_l075_n_93, ZN => VGA_l075_n_119);
  VGA_l075_g12520 : AOI211D0BWP7T port map(A1 => VGA_l075_n_55, A2 => VGA_l075_n_24, B => VGA_l075_n_93, C => VGA_l075_n_78, ZN => VGA_l075_n_118);
  VGA_l075_g12521 : OAI221D0BWP7T port map(A1 => VGA_l075_n_62, A2 => VGA_l075_n_0, B1 => VGA_l075_n_29, B2 => VGA_l075_n_64, C => VGA_l075_n_92, ZN => VGA_l075_n_117);
  VGA_l075_g12522 : OA21D0BWP7T port map(A1 => VGA_l075_n_62, A2 => VGA_l075_n_64, B => VGA_l075_n_92, Z => VGA_l075_n_131);
  VGA_l075_g12523 : AOI22D0BWP7T port map(A1 => VGA_l075_n_66, A2 => VGA_l075_n_31, B1 => VGA_l075_n_47, B2 => VGA_x(2), ZN => VGA_l075_n_129);
  VGA_l075_g12524 : NR3D0BWP7T port map(A1 => VGA_l075_n_80, A2 => VGA_l075_n_73, A3 => VGA_l075_n_61, ZN => VGA_l075_n_128);
  VGA_l075_g12525 : IND2D0BWP7T port map(A1 => VGA_l075_n_37, B1 => VGA_l075_n_102, ZN => VGA_l075_n_127);
  VGA_l075_g12526 : OAI22D0BWP7T port map(A1 => VGA_l075_n_66, A2 => VGA_l075_n_31, B1 => VGA_l075_n_47, B2 => VGA_x(2), ZN => VGA_l075_n_125);
  VGA_l075_g12527 : AN3D0BWP7T port map(A1 => VGA_l075_n_68, A2 => VGA_l075_n_75, A3 => VGA_l075_n_69, Z => VGA_l075_n_124);
  VGA_l075_g12528 : AN2D1BWP7T port map(A1 => VGA_l075_n_88, A2 => VGA_l075_n_68, Z => VGA_l075_n_123);
  VGA_l075_g12529 : AN2D1BWP7T port map(A1 => VGA_l075_n_89, A2 => VGA_l075_n_58, Z => VGA_l075_n_122);
  VGA_l075_g12530 : AOI221D0BWP7T port map(A1 => VGA_l075_n_61, A2 => VGA_draw_count9(0), B1 => VGA_l075_n_56, B2 => VGA_l075_n_25, C => VGA_l075_n_80, ZN => VGA_l075_n_112);
  VGA_l075_g12531 : AO222D0BWP7T port map(A1 => VGA_l075_n_61, A2 => VGA_l075_n_24, B1 => VGA_l075_n_55, B2 => VGA_l075_n_13, C1 => VGA_l075_n_53, C2 => VGA_l075_n_27, Z => VGA_l075_n_111);
  VGA_l075_g12532 : OAI22D0BWP7T port map(A1 => VGA_l075_n_45, A2 => VGA_l075_n_26, B1 => VGA_l075_n_46, B2 => VGA_l075_n_16, ZN => VGA_l075_n_110);
  VGA_l075_g12533 : MAOI22D0BWP7T port map(A1 => VGA_l075_n_50, A2 => VGA_l075_n_35, B1 => VGA_l075_n_50, B2 => VGA_l075_n_35, ZN => VGA_l075_n_109);
  VGA_l075_g12534 : OAI22D0BWP7T port map(A1 => VGA_l075_n_65, A2 => VGA_l075_n_15, B1 => VGA_l075_n_36, B2 => VGA_y(9), ZN => VGA_l075_n_108);
  VGA_l075_g12535 : AOI22D0BWP7T port map(A1 => VGA_l075_n_65, A2 => VGA_l075_n_15, B1 => VGA_l075_n_36, B2 => VGA_y(9), ZN => VGA_l075_n_107);
  VGA_l075_g12536 : MAOI22D0BWP7T port map(A1 => VGA_l075_n_48, A2 => VGA_l075_n_28, B1 => VGA_l075_n_48, B2 => VGA_l075_n_28, ZN => VGA_l075_n_106);
  VGA_l075_g12538 : MAOI22D0BWP7T port map(A1 => VGA_l075_n_38, A2 => VGA_l075_n_19, B1 => VGA_l075_n_38, B2 => VGA_l075_n_19, ZN => VGA_l075_n_116);
  VGA_l075_g12540 : MOAI22D0BWP7T port map(A1 => VGA_l075_n_38, A2 => VGA_l075_n_22, B1 => VGA_l075_n_38, B2 => VGA_l075_n_22, ZN => VGA_l075_n_115);
  VGA_l075_g12541 : MAOI22D0BWP7T port map(A1 => VGA_l075_n_37, A2 => VGA_l075_n_33, B1 => VGA_l075_n_37, B2 => VGA_l075_n_33, ZN => VGA_l075_n_114);
  VGA_l075_g12542 : MOAI22D0BWP7T port map(A1 => VGA_l075_n_37, A2 => VGA_l075_n_23, B1 => VGA_l075_n_37, B2 => VGA_l075_n_23, ZN => VGA_l075_n_113);
  VGA_l075_g12543 : AOI21D0BWP7T port map(A1 => VGA_l075_n_56, A2 => VGA_l075_n_24, B => VGA_l075_n_63, ZN => VGA_l075_n_99);
  VGA_l075_g12544 : NR2D0BWP7T port map(A1 => VGA_l075_n_44, A2 => VGA_l075_n_34, ZN => VGA_l075_n_98);
  VGA_l075_g12545 : IND2D0BWP7T port map(A1 => VGA_l075_n_46, B1 => x_pos_e5(5), ZN => VGA_l075_n_97);
  VGA_l075_g12546 : ND2D0BWP7T port map(A1 => VGA_l075_n_46, A2 => VGA_l075_n_16, ZN => VGA_l075_n_105);
  VGA_l075_g12547 : NR2D0BWP7T port map(A1 => VGA_l075_n_66, A2 => VGA_l075_n_31, ZN => VGA_l075_n_96);
  VGA_l075_g12548 : NR2D0BWP7T port map(A1 => VGA_l075_n_71, A2 => VGA_l075_n_41, ZN => VGA_l075_n_104);
  VGA_l075_g12550 : NR2D0BWP7T port map(A1 => VGA_l075_n_79, A2 => VGA_l075_n_78, ZN => VGA_l075_n_103);
  VGA_l075_g12551 : NR2D0BWP7T port map(A1 => VGA_l075_n_71, A2 => VGA_l075_n_82, ZN => VGA_l075_n_102);
  VGA_l075_g12552 : ND2D0BWP7T port map(A1 => VGA_l075_n_82, A2 => VGA_y(1), ZN => VGA_l075_n_101);
  VGA_l075_g12553 : IND2D0BWP7T port map(A1 => VGA_y(1), B1 => VGA_l075_n_41, ZN => VGA_l075_n_100);
  VGA_l075_g12554 : CKND1BWP7T port map(I => VGA_l075_n_90, ZN => VGA_l075_n_91);
  VGA_l075_g12555 : AOI21D0BWP7T port map(A1 => VGA_l075_n_59, A2 => VGA_l075_n_25, B => VGA_l075_n_73, ZN => VGA_l075_n_86);
  VGA_l075_g12556 : OAI21D0BWP7T port map(A1 => VGA_l075_n_56, A2 => VGA_l075_n_53, B => VGA_l075_n_24, ZN => VGA_l075_n_85);
  VGA_l075_g12557 : AO21D0BWP7T port map(A1 => VGA_l075_n_60, A2 => VGA_l075_n_54, B => VGA_l075_n_62, Z => VGA_l075_n_84);
  VGA_l075_g12558 : IAO21D0BWP7T port map(A1 => VGA_l075_n_60, A2 => VGA_l075_n_13, B => VGA_l075_n_55, ZN => VGA_l075_n_94);
  VGA_l075_g12559 : OAI21D0BWP7T port map(A1 => VGA_l075_n_52, A2 => VGA_draw_count9(1), B => VGA_l075_n_70, ZN => VGA_l075_n_93);
  VGA_l075_g12560 : AOI22D0BWP7T port map(A1 => VGA_l075_n_51, A2 => VGA_x(0), B1 => VGA_x(1), B2 => VGA_l075_n_6, ZN => VGA_l075_n_83);
  VGA_l075_g12561 : OA22D0BWP7T port map(A1 => VGA_l075_n_64, A2 => VGA_l075_n_12, B1 => VGA_l075_n_25, B2 => VGA_l075_n_0, Z => VGA_l075_n_92);
  VGA_l075_g12562 : OAI21D0BWP7T port map(A1 => VGA_l075_n_57, A2 => VGA_l075_n_13, B => VGA_l075_n_69, ZN => VGA_l075_n_90);
  VGA_l075_g12563 : AOI22D0BWP7T port map(A1 => VGA_l075_n_56, A2 => VGA_l075_n_13, B1 => VGA_l075_n_59, B2 => VGA_l075_n_24, ZN => VGA_l075_n_89);
  VGA_l075_g12564 : IAO21D0BWP7T port map(A1 => VGA_l075_n_0, A2 => VGA_l075_n_24, B => VGA_l075_n_79, ZN => VGA_l075_n_88);
  VGA_l075_g12565 : MOAI22D0BWP7T port map(A1 => VGA_l075_n_43, A2 => VGA_y(0), B1 => VGA_l075_n_43, B2 => VGA_y(0), ZN => VGA_l075_n_87);
  VGA_l075_g12568 : INVD0BWP7T port map(I => VGA_l075_n_41, ZN => VGA_l075_n_82);
  VGA_l075_g12569 : CKND1BWP7T port map(I => VGA_l075_n_26, ZN => VGA_l075_n_81);
  VGA_l075_g12570 : NR2D0BWP7T port map(A1 => VGA_l075_n_54, A2 => VGA_draw_count9(1), ZN => VGA_l075_n_80);
  VGA_l075_g12571 : INR2D0BWP7T port map(A1 => VGA_l075_n_63, B1 => VGA_l075_n_25, ZN => VGA_l075_n_79);
  VGA_l075_g12572 : NR2D0BWP7T port map(A1 => VGA_l075_n_0, A2 => VGA_draw_count9(1), ZN => VGA_l075_n_78);
  VGA_l075_g12573 : NR2D0BWP7T port map(A1 => VGA_l075_n_57, A2 => VGA_l075_n_29, ZN => VGA_l075_n_77);
  VGA_l075_g12574 : ND2D0BWP7T port map(A1 => VGA_l075_n_55, A2 => VGA_draw_count9(1), ZN => VGA_l075_n_76);
  VGA_l075_g12575 : ND2D0BWP7T port map(A1 => VGA_l075_n_53, A2 => VGA_l075_n_13, ZN => VGA_l075_n_75);
  VGA_l075_g12576 : ND2D0BWP7T port map(A1 => VGA_l075_n_53, A2 => VGA_draw_count9(1), ZN => VGA_l075_n_74);
  VGA_l075_g12577 : NR2D0BWP7T port map(A1 => VGA_l075_n_56, A2 => VGA_l075_n_59, ZN => VGA_l075_n_67);
  VGA_l075_g12578 : AN2D1BWP7T port map(A1 => VGA_l075_n_63, A2 => VGA_l075_n_27, Z => VGA_l075_n_73);
  VGA_l075_g12579 : NR2D0BWP7T port map(A1 => VGA_l075_n_52, A2 => VGA_l075_n_13, ZN => VGA_l075_n_72);
  VGA_l075_g12580 : ND2D0BWP7T port map(A1 => VGA_l075_n_40, A2 => VGA_l075_n_43, ZN => VGA_l075_n_71);
  VGA_l075_g12581 : IND2D0BWP7T port map(A1 => VGA_l075_n_62, B1 => VGA_l075_n_56, ZN => VGA_l075_n_70);
  VGA_l075_g12582 : ND2D0BWP7T port map(A1 => VGA_l075_n_63, A2 => VGA_l075_n_13, ZN => VGA_l075_n_69);
  VGA_l075_g12583 : IND2D0BWP7T port map(A1 => VGA_l075_n_62, B1 => VGA_l075_n_63, ZN => VGA_l075_n_68);
  VGA_l075_g12584 : INVD0BWP7T port map(I => VGA_l075_n_61, ZN => VGA_l075_n_60);
  VGA_l075_g12585 : INVD0BWP7T port map(I => VGA_l075_n_59, ZN => VGA_l075_n_58);
  VGA_l075_g12586 : INVD1BWP7T port map(I => VGA_l075_n_57, ZN => VGA_l075_n_56);
  VGA_l075_g12587 : INVD0BWP7T port map(I => VGA_l075_n_55, ZN => VGA_l075_n_54);
  VGA_l075_g12588 : INVD0BWP7T port map(I => VGA_l075_n_53, ZN => VGA_l075_n_52);
  VGA_l075_g12589 : IAO21D0BWP7T port map(A1 => VGA_x(1), A2 => VGA_l075_n_6, B => x_pos_e5(0), ZN => VGA_l075_n_51);
  VGA_l075_g12590 : OAI21D0BWP7T port map(A1 => VGA_l075_n_7, A2 => x_pos_e5(4), B => VGA_l075_n_26, ZN => VGA_l075_n_66);
  VGA_l075_g12591 : AOI21D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l075_n_5, B => VGA_l075_n_28, ZN => VGA_l075_n_65);
  VGA_l075_g12592 : IND2D0BWP7T port map(A1 => VGA_l075_n_30, B1 => VGA_draw_count9(4), ZN => VGA_l075_n_64);
  VGA_l075_g12593 : INR2D0BWP7T port map(A1 => VGA_draw_count9(4), B1 => VGA_l075_n_17, ZN => VGA_l075_n_63);
  VGA_l075_g12594 : INR2D0BWP7T port map(A1 => VGA_l075_n_29, B1 => VGA_l075_n_27, ZN => VGA_l075_n_62);
  VGA_l075_g12596 : NR2D0BWP7T port map(A1 => VGA_l075_n_14, A2 => VGA_draw_count9(4), ZN => VGA_l075_n_61);
  VGA_l075_g12597 : NR2D0BWP7T port map(A1 => VGA_l075_n_30, A2 => VGA_draw_count9(4), ZN => VGA_l075_n_59);
  VGA_l075_g12598 : IND2D0BWP7T port map(A1 => VGA_l075_n_14, B1 => VGA_draw_count9(4), ZN => VGA_l075_n_57);
  VGA_l075_g12599 : NR2D0BWP7T port map(A1 => VGA_l075_n_17, A2 => VGA_draw_count9(4), ZN => VGA_l075_n_55);
  VGA_l075_g12600 : NR2D0BWP7T port map(A1 => VGA_l075_n_18, A2 => VGA_draw_count9(4), ZN => VGA_l075_n_53);
  VGA_l075_g12601 : CKND1BWP7T port map(I => VGA_l075_n_43, ZN => VGA_l075_n_42);
  VGA_l075_g12602 : CKND1BWP7T port map(I => VGA_l075_n_40, ZN => VGA_l075_n_39);
  VGA_l075_g12603 : MOAI22D0BWP7T port map(A1 => VGA_y(8), A2 => y_pos_e5(8), B1 => VGA_y(8), B2 => y_pos_e5(8), ZN => VGA_l075_n_50);
  VGA_l075_g12604 : MOAI22D0BWP7T port map(A1 => VGA_x(7), A2 => x_pos_e5(7), B1 => VGA_x(7), B2 => x_pos_e5(7), ZN => VGA_l075_n_49);
  VGA_l075_g12605 : MOAI22D0BWP7T port map(A1 => VGA_y(7), A2 => y_pos_e5(7), B1 => VGA_y(7), B2 => y_pos_e5(7), ZN => VGA_l075_n_48);
  VGA_l075_g12606 : MAOI22D0BWP7T port map(A1 => VGA_x(3), A2 => x_pos_e5(3), B1 => VGA_x(3), B2 => x_pos_e5(3), ZN => VGA_l075_n_47);
  VGA_l075_g12607 : MOAI22D0BWP7T port map(A1 => VGA_x(6), A2 => x_pos_e5(6), B1 => VGA_x(6), B2 => x_pos_e5(6), ZN => VGA_l075_n_46);
  VGA_l075_g12608 : MOAI22D0BWP7T port map(A1 => VGA_x(5), A2 => x_pos_e5(5), B1 => VGA_x(5), B2 => x_pos_e5(5), ZN => VGA_l075_n_45);
  VGA_l075_g12609 : MAOI22D0BWP7T port map(A1 => VGA_y(5), A2 => y_pos_e5(5), B1 => VGA_y(5), B2 => y_pos_e5(5), ZN => VGA_l075_n_44);
  VGA_l075_g12610 : MOAI22D0BWP7T port map(A1 => VGA_y(1), A2 => y_pos_e5(1), B1 => VGA_y(1), B2 => y_pos_e5(1), ZN => VGA_l075_n_43);
  VGA_l075_g12611 : MOAI22D0BWP7T port map(A1 => VGA_y(2), A2 => y_pos_e5(2), B1 => VGA_y(2), B2 => y_pos_e5(2), ZN => VGA_l075_n_41);
  VGA_l075_g12612 : MOAI22D0BWP7T port map(A1 => VGA_y(0), A2 => y_pos_e5(0), B1 => VGA_y(0), B2 => y_pos_e5(0), ZN => VGA_l075_n_40);
  VGA_l075_g12613 : MAOI22D0BWP7T port map(A1 => VGA_y(4), A2 => y_pos_e5(4), B1 => VGA_y(4), B2 => y_pos_e5(4), ZN => VGA_l075_n_38);
  VGA_l075_g12614 : MOAI22D0BWP7T port map(A1 => VGA_y(3), A2 => y_pos_e5(3), B1 => VGA_y(3), B2 => y_pos_e5(3), ZN => VGA_l075_n_37);
  VGA_l075_g12615 : INVD1BWP7T port map(I => VGA_l075_n_25, ZN => VGA_l075_n_24);
  VGA_l075_g12616 : IND2D0BWP7T port map(A1 => VGA_y(8), B1 => y_pos_e5(8), ZN => VGA_l075_n_36);
  VGA_l075_g12617 : INR2D0BWP7T port map(A1 => y_pos_e5(7), B1 => VGA_y(7), ZN => VGA_l075_n_35);
  VGA_l075_g12618 : IND2D0BWP7T port map(A1 => y_pos_e5(4), B1 => VGA_y(4), ZN => VGA_l075_n_34);
  VGA_l075_g12619 : IND2D0BWP7T port map(A1 => y_pos_e5(2), B1 => VGA_y(2), ZN => VGA_l075_n_33);
  VGA_l075_g12620 : IND2D0BWP7T port map(A1 => x_pos_e5(6), B1 => VGA_x(6), ZN => VGA_l075_n_32);
  VGA_l075_g12621 : IND2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_e5(3), ZN => VGA_l075_n_31);
  VGA_l075_g12622 : ND2D0BWP7T port map(A1 => VGA_draw_count9(2), A2 => VGA_draw_count9(3), ZN => VGA_l075_n_30);
  VGA_l075_g12623 : ND2D0BWP7T port map(A1 => VGA_l075_n_3, A2 => VGA_draw_count9(0), ZN => VGA_l075_n_29);
  VGA_l075_g12624 : NR2D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l075_n_5, ZN => VGA_l075_n_28);
  VGA_l075_g12625 : NR2D0BWP7T port map(A1 => VGA_l075_n_3, A2 => VGA_draw_count9(0), ZN => VGA_l075_n_27);
  VGA_l075_g12626 : ND2D0BWP7T port map(A1 => VGA_l075_n_7, A2 => x_pos_e5(4), ZN => VGA_l075_n_26);
  VGA_l075_g12627 : ND2D0BWP7T port map(A1 => VGA_draw_count9(1), A2 => VGA_draw_count9(0), ZN => VGA_l075_n_25);
  VGA_l075_g12629 : CKND1BWP7T port map(I => VGA_l075_n_13, ZN => VGA_l075_n_12);
  VGA_l075_g12630 : IND2D0BWP7T port map(A1 => VGA_y(4), B1 => y_pos_e5(4), ZN => VGA_l075_n_11);
  VGA_l075_g12631 : ND2D0BWP7T port map(A1 => VGA_l075_n_8, A2 => y_pos_e5(2), ZN => VGA_l075_n_23);
  VGA_l075_g12632 : NR2D0BWP7T port map(A1 => VGA_l075_n_9, A2 => y_pos_e5(3), ZN => VGA_l075_n_22);
  VGA_l075_g12633 : INR2D0BWP7T port map(A1 => x_pos_e5(7), B1 => VGA_x(7), ZN => VGA_l075_n_21);
  VGA_l075_g12634 : ND2D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l075_n_10, ZN => VGA_l075_n_20);
  VGA_l075_g12635 : INR2D0BWP7T port map(A1 => y_pos_e5(3), B1 => VGA_y(3), ZN => VGA_l075_n_19);
  VGA_l075_g12636 : IND2D0BWP7T port map(A1 => VGA_draw_count9(2), B1 => VGA_draw_count9(3), ZN => VGA_l075_n_18);
  VGA_l075_g12637 : IND2D0BWP7T port map(A1 => VGA_draw_count9(3), B1 => VGA_draw_count9(2), ZN => VGA_l075_n_17);
  VGA_l075_g12638 : INR2D0BWP7T port map(A1 => VGA_x(5), B1 => x_pos_e5(5), ZN => VGA_l075_n_16);
  VGA_l075_g12639 : IND2D0BWP7T port map(A1 => y_pos_e5(5), B1 => VGA_y(5), ZN => VGA_l075_n_15);
  VGA_l075_g12640 : OR2D0BWP7T port map(A1 => VGA_draw_count9(2), A2 => VGA_draw_count9(3), Z => VGA_l075_n_14);
  VGA_l075_g12641 : NR2D0BWP7T port map(A1 => VGA_draw_count9(1), A2 => VGA_draw_count9(0), ZN => VGA_l075_n_13);
  VGA_l075_g12642 : CKND1BWP7T port map(I => x_pos_e5(8), ZN => VGA_l075_n_10);
  VGA_l075_g12643 : CKND1BWP7T port map(I => VGA_y(3), ZN => VGA_l075_n_9);
  VGA_l075_g12644 : CKND1BWP7T port map(I => VGA_y(2), ZN => VGA_l075_n_8);
  VGA_l075_g12645 : CKND1BWP7T port map(I => VGA_x(4), ZN => VGA_l075_n_7);
  VGA_l075_g12646 : CKND1BWP7T port map(I => x_pos_e5(1), ZN => VGA_l075_n_6);
  VGA_l075_g12647 : CKND1BWP7T port map(I => y_pos_e5(6), ZN => VGA_l075_n_5);
  VGA_l075_g12648 : CKND1BWP7T port map(I => y_pos_e5(1), ZN => VGA_l075_n_4);
  VGA_l075_g12649 : INVD0BWP7T port map(I => VGA_draw_count9(1), ZN => VGA_l075_n_3);
  VGA_l075_g2 : MUX2ND0BWP7T port map(I0 => VGA_y(3), I1 => VGA_l075_n_9, S => VGA_l075_n_38, ZN => VGA_l075_n_2);
  VGA_l075_g12650 : MUX2ND0BWP7T port map(I0 => VGA_l075_n_8, I1 => VGA_y(2), S => VGA_l075_n_37, ZN => VGA_l075_n_1);
  VGA_l075_g12651 : IND2D1BWP7T port map(A1 => VGA_l075_n_18, B1 => VGA_draw_count9(4), ZN => VGA_l075_n_0);
  VGA_l075_g12652 : INVD0BWP7T port map(I => VGA_l075_n_66, ZN => VGA_l075_n_95);
  VGA_l076_g12402 : OAI211D0BWP7T port map(A1 => VGA_l076_n_76, A2 => VGA_l076_n_195, B => VGA_l076_n_243, C => VGA_l076_n_223, ZN => VGA_r10);
  VGA_l076_g12403 : AOI211D0BWP7T port map(A1 => VGA_l076_n_206, A2 => VGA_l076_n_111, B => VGA_l076_n_242, C => VGA_l076_n_225, ZN => VGA_l076_n_243);
  VGA_l076_g12404 : OAI211D0BWP7T port map(A1 => VGA_l076_n_162, A2 => VGA_l076_n_216, B => VGA_l076_n_241, C => VGA_l076_n_238, ZN => VGA_l076_n_242);
  VGA_l076_g12405 : NR4D0BWP7T port map(A1 => VGA_l076_n_239, A2 => VGA_l076_n_227, A3 => VGA_l076_n_219, A4 => VGA_l076_n_220, ZN => VGA_l076_n_241);
  VGA_l076_g12406 : OAI211D0BWP7T port map(A1 => VGA_l076_n_91, A2 => VGA_l076_n_212, B => VGA_l076_n_237, C => VGA_l076_n_235, ZN => VGA_g10);
  VGA_l076_g12407 : NR4D0BWP7T port map(A1 => VGA_l076_n_233, A2 => VGA_l076_n_191, A3 => VGA_l076_n_151, A4 => VGA_l076_n_138, ZN => VGA_l076_n_239);
  VGA_l076_g12408 : NR4D0BWP7T port map(A1 => VGA_l076_n_226, A2 => VGA_l076_n_228, A3 => VGA_l076_n_221, A4 => VGA_l076_n_192, ZN => VGA_l076_n_238);
  VGA_l076_g12409 : AOI211D0BWP7T port map(A1 => VGA_l076_n_206, A2 => VGA_l076_n_117, B => VGA_l076_n_236, C => VGA_l076_n_218, ZN => VGA_l076_n_237);
  VGA_l076_g12410 : OAI211D0BWP7T port map(A1 => VGA_l076_n_99, A2 => VGA_l076_n_195, B => VGA_l076_n_230, C => VGA_l076_n_224, ZN => VGA_l076_n_236);
  VGA_l076_g12411 : AOI211D0BWP7T port map(A1 => VGA_l076_n_211, A2 => VGA_l076_n_137, B => VGA_l076_n_231, C => VGA_l076_n_213, ZN => VGA_l076_n_235);
  VGA_l076_g12412 : OAI32D0BWP7T port map(A1 => VGA_l076_n_24, A2 => VGA_l076_n_60, A3 => VGA_l076_n_216, B1 => VGA_l076_n_94, B2 => VGA_l076_n_215, ZN => VGA_b10);
  VGA_l076_g12413 : ND4D0BWP7T port map(A1 => VGA_l076_n_210, A2 => VGA_l076_n_189, A3 => VGA_l076_n_176, A4 => VGA_l076_n_165, ZN => VGA_l076_n_233);
  VGA_l076_g12414 : OAI211D0BWP7T port map(A1 => VGA_l076_n_191, A2 => VGA_l076_n_209, B => VGA_l076_n_204, C => VGA_l076_n_199, ZN => VGA_enable10);
  VGA_l076_g12415 : OAI22D0BWP7T port map(A1 => VGA_l076_n_217, A2 => VGA_l076_n_139, B1 => VGA_l076_n_207, B2 => VGA_l076_n_131, ZN => VGA_l076_n_231);
  VGA_l076_g12416 : AOI31D0BWP7T port map(A1 => VGA_l076_n_190, A2 => VGA_l076_n_182, A3 => VGA_l076_n_77, B => VGA_l076_n_229, ZN => VGA_l076_n_230);
  VGA_l076_g12417 : AOI21D0BWP7T port map(A1 => VGA_l076_n_103, A2 => VGA_l076_n_86, B => VGA_l076_n_216, ZN => VGA_l076_n_229);
  VGA_l076_g12418 : AOI31D0BWP7T port map(A1 => VGA_l076_n_145, A2 => VGA_l076_n_88, A3 => VGA_l076_n_75, B => VGA_l076_n_217, ZN => VGA_l076_n_228);
  VGA_l076_g12419 : AOI31D0BWP7T port map(A1 => VGA_l076_n_122, A2 => VGA_l076_n_118, A3 => VGA_l076_n_60, B => VGA_l076_n_214, ZN => VGA_l076_n_227);
  VGA_l076_g12420 : AOI31D0BWP7T port map(A1 => VGA_l076_n_142, A2 => VGA_l076_n_122, A3 => VGA_l076_n_88, B => VGA_l076_n_215, ZN => VGA_l076_n_226);
  VGA_l076_g12421 : AOI22D0BWP7T port map(A1 => VGA_l076_n_205, A2 => VGA_l076_n_195, B1 => VGA_l076_n_119, B2 => VGA_l076_n_89, ZN => VGA_l076_n_225);
  VGA_l076_g12422 : AO21D0BWP7T port map(A1 => VGA_l076_n_123, A2 => VGA_l076_n_91, B => VGA_l076_n_215, Z => VGA_l076_n_224);
  VGA_l076_g12423 : OA21D0BWP7T port map(A1 => VGA_l076_n_208, A2 => VGA_l076_n_157, B => VGA_l076_n_222, Z => VGA_l076_n_223);
  VGA_l076_g12424 : AO31D0BWP7T port map(A1 => VGA_l076_n_135, A2 => VGA_l076_n_68, A3 => VGA_l076_n_69, B => VGA_l076_n_204, Z => VGA_l076_n_222);
  VGA_l076_g12425 : AOI21D0BWP7T port map(A1 => VGA_l076_n_89, A2 => VGA_l076_n_52, B => VGA_l076_n_212, ZN => VGA_l076_n_221);
  VGA_l076_g12426 : AOI31D0BWP7T port map(A1 => VGA_l076_n_132, A2 => VGA_l076_n_76, A3 => VGA_l076_n_58, B => VGA_l076_n_207, ZN => VGA_l076_n_220);
  VGA_l076_g12427 : OA21D0BWP7T port map(A1 => VGA_l076_n_134, A2 => VGA_l076_n_90, B => VGA_l076_n_211, Z => VGA_l076_n_219);
  VGA_l076_g12428 : AOI21D0BWP7T port map(A1 => VGA_l076_n_88, A2 => VGA_l076_n_0, B => VGA_l076_n_204, ZN => VGA_l076_n_218);
  VGA_l076_g12429 : AOI32D0BWP7T port map(A1 => VGA_l076_n_190, A2 => VGA_l076_n_181, A3 => VGA_l076_n_38, B1 => VGA_l076_n_202, B2 => VGA_l076_n_154, ZN => VGA_l076_n_214);
  VGA_l076_g12430 : AOI21D0BWP7T port map(A1 => VGA_l076_n_103, A2 => VGA_l076_n_68, B => VGA_l076_n_208, ZN => VGA_l076_n_213);
  VGA_l076_g12431 : AOI22D0BWP7T port map(A1 => VGA_l076_n_203, A2 => VGA_l076_n_156, B1 => VGA_l076_n_202, B2 => VGA_l076_n_143, ZN => VGA_l076_n_217);
  VGA_l076_g12432 : AOI22D0BWP7T port map(A1 => VGA_l076_n_202, A2 => VGA_l076_n_160, B1 => VGA_l076_n_203, B2 => VGA_l076_n_144, ZN => VGA_l076_n_216);
  VGA_l076_g12433 : AOI32D0BWP7T port map(A1 => VGA_l076_n_198, A2 => VGA_l076_n_1, A3 => VGA_l076_n_104, B1 => VGA_l076_n_203, B2 => VGA_l076_n_155, ZN => VGA_l076_n_215);
  VGA_l076_g12434 : OAI31D0BWP7T port map(A1 => VGA_l076_n_2, A2 => VGA_l076_n_127, A3 => VGA_l076_n_179, B => VGA_l076_n_201, ZN => VGA_l076_n_210);
  VGA_l076_g12435 : NR4D0BWP7T port map(A1 => VGA_l076_n_200, A2 => VGA_l076_n_186, A3 => VGA_l076_n_182, A4 => VGA_l076_n_185, ZN => VGA_l076_n_209);
  VGA_l076_g12436 : MAOI22D0BWP7T port map(A1 => VGA_l076_n_196, A2 => VGA_l076_n_170, B1 => VGA_l076_n_191, B2 => VGA_l076_n_165, ZN => VGA_l076_n_212);
  VGA_l076_g12437 : OAI22D0BWP7T port map(A1 => VGA_l076_n_197, A2 => VGA_l076_n_171, B1 => VGA_l076_n_193, B2 => VGA_l076_n_150, ZN => VGA_l076_n_211);
  VGA_l076_g12438 : CKND1BWP7T port map(I => VGA_l076_n_206, ZN => VGA_l076_n_205);
  VGA_l076_g12439 : AOI22D0BWP7T port map(A1 => VGA_l076_n_196, A2 => VGA_l076_n_169, B1 => VGA_l076_n_194, B2 => VGA_l076_n_151, ZN => VGA_l076_n_208);
  VGA_l076_g12440 : MAOI22D0BWP7T port map(A1 => VGA_l076_n_196, A2 => VGA_l076_n_151, B1 => VGA_l076_n_193, B2 => VGA_l076_n_168, ZN => VGA_l076_n_207);
  VGA_l076_g12441 : OAI22D0BWP7T port map(A1 => VGA_l076_n_197, A2 => VGA_l076_n_167, B1 => VGA_l076_n_191, B2 => VGA_l076_n_176, ZN => VGA_l076_n_206);
  VGA_l076_g12442 : MAOI22D0BWP7T port map(A1 => VGA_l076_n_196, A2 => VGA_l076_n_140, B1 => VGA_l076_n_193, B2 => VGA_l076_n_167, ZN => VGA_l076_n_204);
  VGA_l076_g12443 : INR2D0BWP7T port map(A1 => VGA_l076_n_198, B1 => VGA_l076_n_114, ZN => VGA_l076_n_203);
  VGA_l076_g12444 : INR2D0BWP7T port map(A1 => VGA_l076_n_198, B1 => VGA_l076_n_113, ZN => VGA_l076_n_202);
  VGA_l076_g12445 : CKND1BWP7T port map(I => VGA_l076_n_200, ZN => VGA_l076_n_201);
  VGA_l076_g12446 : OAI21D0BWP7T port map(A1 => VGA_l076_n_177, A2 => VGA_l076_n_161, B => VGA_l076_n_194, ZN => VGA_l076_n_199);
  VGA_l076_g12447 : ND3D0BWP7T port map(A1 => VGA_l076_n_188, A2 => VGA_l076_n_176, A3 => VGA_l076_n_165, ZN => VGA_l076_n_200);
  VGA_l076_g12448 : INVD0BWP7T port map(I => VGA_l076_n_197, ZN => VGA_l076_n_196);
  VGA_l076_g12449 : INR2D0BWP7T port map(A1 => VGA_l076_n_185, B1 => VGA_l076_n_191, ZN => VGA_l076_n_198);
  VGA_l076_g12450 : ND2D0BWP7T port map(A1 => VGA_l076_n_190, A2 => VGA_l076_n_184, ZN => VGA_l076_n_197);
  VGA_l076_g12451 : CKND1BWP7T port map(I => VGA_l076_n_193, ZN => VGA_l076_n_194);
  VGA_l076_g12452 : AOI211D0BWP7T port map(A1 => VGA_l076_n_122, A2 => VGA_l076_n_74, B => VGA_l076_n_191, C => VGA_l076_n_183, ZN => VGA_l076_n_192);
  VGA_l076_g12453 : IND2D0BWP7T port map(A1 => VGA_l076_n_189, B1 => VGA_l076_n_190, ZN => VGA_l076_n_195);
  VGA_l076_g12454 : ND2D0BWP7T port map(A1 => VGA_l076_n_190, A2 => VGA_l076_n_164, ZN => VGA_l076_n_193);
  VGA_l076_g12455 : INVD1BWP7T port map(I => VGA_l076_n_191, ZN => VGA_l076_n_190);
  VGA_l076_g12456 : OAI221D0BWP7T port map(A1 => VGA_l076_n_49, A2 => VGA_l076_n_32, B1 => VGA_l076_n_20, B2 => VGA_l076_n_21, C => VGA_l076_n_187, ZN => VGA_l076_n_191);
  VGA_l076_g12457 : AOI22D0BWP7T port map(A1 => VGA_l076_n_184, A2 => VGA_l076_n_161, B1 => VGA_l076_n_170, B2 => VGA_l076_n_164, ZN => VGA_l076_n_188);
  VGA_l076_g12458 : AOI33D0BWP7T port map(A1 => VGA_l076_n_184, A2 => VGA_l076_n_143, A3 => VGA_l076_n_113, B1 => VGA_l076_n_164, B2 => VGA_l076_n_156, B3 => VGA_l076_n_114, ZN => VGA_l076_n_189);
  VGA_l076_g12459 : AOI211D0BWP7T port map(A1 => VGA_l076_n_173, A2 => VGA_l076_n_136, B => VGA_l076_n_178, C => VGA_l076_n_120, ZN => VGA_l076_n_187);
  VGA_l076_g12460 : OA21D0BWP7T port map(A1 => VGA_l076_n_180, A2 => VGA_l076_n_170, B => VGA_l076_n_184, Z => VGA_l076_n_186);
  VGA_l076_g12461 : NR2D0BWP7T port map(A1 => VGA_l076_n_179, A2 => VGA_l076_n_115, ZN => VGA_l076_n_185);
  VGA_l076_g12462 : NR2D0BWP7T port map(A1 => VGA_l076_n_179, A2 => VGA_l076_n_116, ZN => VGA_l076_n_184);
  VGA_l076_g12463 : CKND1BWP7T port map(I => VGA_l076_n_182, ZN => VGA_l076_n_183);
  VGA_l076_g12464 : AO32D0BWP7T port map(A1 => VGA_l076_n_166, A2 => VGA_l076_n_102, A3 => VGA_l076_n_37, B1 => VGA_l076_n_175, B2 => VGA_y(4), Z => VGA_l076_n_181);
  VGA_l076_g12465 : OAI22D0BWP7T port map(A1 => VGA_l076_n_172, A2 => VGA_l076_n_113, B1 => VGA_l076_n_174, B2 => VGA_l076_n_38, ZN => VGA_l076_n_182);
  VGA_l076_g12466 : IND2D0BWP7T port map(A1 => VGA_l076_n_177, B1 => VGA_l076_n_167, ZN => VGA_l076_n_180);
  VGA_l076_g12467 : MOAI22D0BWP7T port map(A1 => VGA_l076_n_163, A2 => VGA_l076_n_136, B1 => VGA_l076_n_21, B2 => VGA_l076_n_20, ZN => VGA_l076_n_178);
  VGA_l076_g12468 : AOI22D0BWP7T port map(A1 => VGA_l076_n_166, A2 => y_pos_e6(4), B1 => VGA_l076_n_159, B2 => VGA_l076_n_11, ZN => VGA_l076_n_179);
  VGA_l076_g12469 : ND2D0BWP7T port map(A1 => VGA_l076_n_168, A2 => VGA_l076_n_171, ZN => VGA_l076_n_177);
  VGA_l076_g12470 : ND2D0BWP7T port map(A1 => VGA_l076_n_164, A2 => VGA_l076_n_140, ZN => VGA_l076_n_176);
  VGA_l076_g12471 : CKND1BWP7T port map(I => VGA_l076_n_174, ZN => VGA_l076_n_175);
  VGA_l076_g12472 : OAI211D0BWP7T port map(A1 => VGA_l076_n_96, A2 => VGA_l076_n_129, B => VGA_l076_n_153, C => VGA_l076_n_105, ZN => VGA_l076_n_173);
  VGA_l076_g12473 : ND3D0BWP7T port map(A1 => VGA_l076_n_154, A2 => VGA_l076_n_158, A3 => VGA_l076_n_115, ZN => VGA_l076_n_172);
  VGA_l076_g12474 : ND3D0BWP7T port map(A1 => VGA_l076_n_159, A2 => VGA_l076_n_102, A3 => VGA_l076_n_37, ZN => VGA_l076_n_174);
  VGA_l076_g12475 : CKND1BWP7T port map(I => VGA_l076_n_168, ZN => VGA_l076_n_169);
  VGA_l076_g12476 : ND2D0BWP7T port map(A1 => VGA_l076_n_156, A2 => VGA_l076_n_114, ZN => VGA_l076_n_171);
  VGA_l076_g12477 : AN2D1BWP7T port map(A1 => VGA_l076_n_154, A2 => VGA_l076_n_113, Z => VGA_l076_n_170);
  VGA_l076_g12478 : ND2D0BWP7T port map(A1 => VGA_l076_n_160, A2 => VGA_l076_n_113, ZN => VGA_l076_n_168);
  VGA_l076_g12479 : ND2D0BWP7T port map(A1 => VGA_l076_n_155, A2 => VGA_l076_n_114, ZN => VGA_l076_n_167);
  VGA_l076_g12480 : AOI221D0BWP7T port map(A1 => VGA_l076_n_125, A2 => VGA_l076_n_95, B1 => VGA_l076_n_45, B2 => VGA_l076_n_81, C => VGA_l076_n_152, ZN => VGA_l076_n_163);
  VGA_l076_g12481 : AN4D1BWP7T port map(A1 => VGA_l076_n_141, A2 => VGA_l076_n_103, A3 => VGA_l076_n_89, A4 => VGA_l076_n_0, Z => VGA_l076_n_162);
  VGA_l076_g12482 : NR3D0BWP7T port map(A1 => VGA_l076_n_149, A2 => VGA_l076_n_44, A3 => VGA_y(4), ZN => VGA_l076_n_166);
  VGA_l076_g12483 : IND3D0BWP7T port map(A1 => VGA_l076_n_127, B1 => VGA_l076_n_2, B2 => VGA_l076_n_158, ZN => VGA_l076_n_165);
  VGA_l076_g12484 : AN2D1BWP7T port map(A1 => VGA_l076_n_158, A2 => VGA_l076_n_116, Z => VGA_l076_n_164);
  VGA_l076_g12485 : IINR4D0BWP7T port map(A1 => VGA_l076_n_122, A2 => VGA_l076_n_69, B1 => VGA_l076_n_133, B2 => VGA_l076_n_77, ZN => VGA_l076_n_157);
  VGA_l076_g12486 : IND2D0BWP7T port map(A1 => VGA_l076_n_151, B1 => VGA_l076_n_150, ZN => VGA_l076_n_161);
  VGA_l076_g12487 : NR3D0BWP7T port map(A1 => VGA_l076_n_148, A2 => VGA_l076_n_87, A3 => VGA_l076_n_40, ZN => VGA_l076_n_160);
  VGA_l076_g12488 : INR2D0BWP7T port map(A1 => VGA_l076_n_44, B1 => VGA_l076_n_149, ZN => VGA_l076_n_159);
  VGA_l076_g12489 : AOI211D0BWP7T port map(A1 => VGA_l076_n_44, A2 => VGA_l076_n_34, B => VGA_l076_n_149, C => VGA_l076_n_98, ZN => VGA_l076_n_158);
  VGA_l076_g12490 : AOI22D0BWP7T port map(A1 => VGA_l076_n_146, A2 => VGA_l076_n_126, B1 => VGA_l076_n_45, B2 => VGA_l076_n_26, ZN => VGA_l076_n_153);
  VGA_l076_g12491 : OAI22D0BWP7T port map(A1 => VGA_l076_n_146, A2 => VGA_l076_n_130, B1 => VGA_l076_n_97, B2 => VGA_x(5), ZN => VGA_l076_n_152);
  VGA_l076_g12492 : INR3D0BWP7T port map(A1 => VGA_l076_n_148, B1 => VGA_l076_n_40, B2 => VGA_l076_n_87, ZN => VGA_l076_n_156);
  VGA_l076_g12493 : AN3D0BWP7T port map(A1 => VGA_l076_n_147, A2 => VGA_l076_n_87, A3 => VGA_l076_n_39, Z => VGA_l076_n_155);
  VGA_l076_g12494 : INR3D0BWP7T port map(A1 => VGA_l076_n_87, B1 => VGA_l076_n_40, B2 => VGA_l076_n_147, ZN => VGA_l076_n_154);
  VGA_l076_g12495 : AN2D1BWP7T port map(A1 => VGA_l076_n_144, A2 => VGA_l076_n_114, Z => VGA_l076_n_151);
  VGA_l076_g12496 : ND2D0BWP7T port map(A1 => VGA_l076_n_143, A2 => VGA_l076_n_113, ZN => VGA_l076_n_150);
  VGA_l076_g12497 : IND4D0BWP7T port map(A1 => VGA_l076_n_108, B1 => VGA_l076_n_109, B2 => VGA_l076_n_106, B3 => VGA_l076_n_107, ZN => VGA_l076_n_149);
  VGA_l076_g12498 : AN3D0BWP7T port map(A1 => VGA_l076_n_128, A2 => VGA_l076_n_70, A3 => VGA_l076_n_76, Z => VGA_l076_n_145);
  VGA_l076_g12499 : OAI221D0BWP7T port map(A1 => VGA_l076_n_101, A2 => y_pos_e6(1), B1 => VGA_l076_n_4, B2 => VGA_l076_n_82, C => VGA_l076_n_100, ZN => VGA_l076_n_148);
  VGA_l076_g12500 : OAI211D0BWP7T port map(A1 => y_pos_e6(1), A2 => VGA_l076_n_41, B => VGA_l076_n_121, C => VGA_l076_n_101, ZN => VGA_l076_n_147);
  VGA_l076_g12501 : MAOI222D0BWP7T port map(A => VGA_x(2), B => x_pos_e6(2), C => VGA_l076_n_83, ZN => VGA_l076_n_146);
  VGA_l076_g12502 : AN3D0BWP7T port map(A1 => VGA_l076_n_124, A2 => VGA_l076_n_94, A3 => VGA_l076_n_92, Z => VGA_l076_n_142);
  VGA_l076_g12503 : INR3D0BWP7T port map(A1 => VGA_l076_n_128, B1 => VGA_l076_n_72, B2 => VGA_l076_n_77, ZN => VGA_l076_n_141);
  VGA_l076_g12504 : AOI211D0BWP7T port map(A1 => VGA_l076_n_101, A2 => VGA_l076_n_100, B => VGA_l076_n_39, C => VGA_l076_n_43, ZN => VGA_l076_n_144);
  VGA_l076_g12505 : AN4D1BWP7T port map(A1 => VGA_l076_n_101, A2 => VGA_l076_n_100, A3 => VGA_l076_n_42, A4 => VGA_l076_n_40, Z => VGA_l076_n_143);
  VGA_l076_g12506 : INR2D0BWP7T port map(A1 => VGA_l076_n_122, B1 => VGA_l076_n_72, ZN => VGA_l076_n_139);
  VGA_l076_g12507 : AN2D1BWP7T port map(A1 => VGA_l076_n_112, A2 => VGA_l076_n_52, Z => VGA_l076_n_138);
  VGA_l076_g12508 : ND2D0BWP7T port map(A1 => VGA_l076_n_123, A2 => VGA_l076_n_131, ZN => VGA_l076_n_137);
  VGA_l076_g12509 : INR2D0BWP7T port map(A1 => VGA_l076_n_104, B1 => VGA_l076_n_1, ZN => VGA_l076_n_140);
  VGA_l076_g12510 : OA221D0BWP7T port map(A1 => VGA_l076_n_67, A2 => VGA_draw_count10(1), B1 => VGA_l076_n_24, B2 => VGA_l076_n_54, C => VGA_l076_n_74, Z => VGA_l076_n_135);
  VGA_l076_g12511 : OAI211D0BWP7T port map(A1 => VGA_draw_count10(1), A2 => VGA_l076_n_58, B => VGA_l076_n_84, C => VGA_l076_n_74, ZN => VGA_l076_n_134);
  VGA_l076_g12512 : OAI211D0BWP7T port map(A1 => VGA_l076_n_13, A2 => VGA_l076_n_54, B => VGA_l076_n_85, C => VGA_l076_n_75, ZN => VGA_l076_n_133);
  VGA_l076_g12513 : OA21D0BWP7T port map(A1 => VGA_l076_n_14, A2 => VGA_l076_n_3, B => VGA_l076_n_124, Z => VGA_l076_n_132);
  VGA_l076_g12514 : ND2D0BWP7T port map(A1 => VGA_l076_n_110, A2 => VGA_l076_n_105, ZN => VGA_l076_n_136);
  VGA_l076_g12515 : CKND1BWP7T port map(I => VGA_l076_n_129, ZN => VGA_l076_n_130);
  VGA_l076_g12516 : CKND1BWP7T port map(I => VGA_l076_n_125, ZN => VGA_l076_n_126);
  VGA_l076_g12517 : IND2D0BWP7T port map(A1 => VGA_l076_n_100, B1 => y_pos_e6(1), ZN => VGA_l076_n_121);
  VGA_l076_g12518 : MOAI22D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l076_n_10, B1 => VGA_l076_n_49, B2 => VGA_l076_n_32, ZN => VGA_l076_n_120);
  VGA_l076_g12519 : AOI21D0BWP7T port map(A1 => VGA_l076_n_59, A2 => VGA_l076_n_27, B => VGA_l076_n_93, ZN => VGA_l076_n_119);
  VGA_l076_g12520 : AOI211D0BWP7T port map(A1 => VGA_l076_n_55, A2 => VGA_l076_n_24, B => VGA_l076_n_93, C => VGA_l076_n_78, ZN => VGA_l076_n_118);
  VGA_l076_g12521 : OAI221D0BWP7T port map(A1 => VGA_l076_n_62, A2 => VGA_l076_n_0, B1 => VGA_l076_n_29, B2 => VGA_l076_n_64, C => VGA_l076_n_92, ZN => VGA_l076_n_117);
  VGA_l076_g12522 : OA21D0BWP7T port map(A1 => VGA_l076_n_62, A2 => VGA_l076_n_64, B => VGA_l076_n_92, Z => VGA_l076_n_131);
  VGA_l076_g12523 : AOI22D0BWP7T port map(A1 => VGA_l076_n_66, A2 => VGA_l076_n_31, B1 => VGA_l076_n_47, B2 => VGA_x(2), ZN => VGA_l076_n_129);
  VGA_l076_g12524 : NR3D0BWP7T port map(A1 => VGA_l076_n_80, A2 => VGA_l076_n_73, A3 => VGA_l076_n_61, ZN => VGA_l076_n_128);
  VGA_l076_g12525 : IND2D0BWP7T port map(A1 => VGA_l076_n_37, B1 => VGA_l076_n_102, ZN => VGA_l076_n_127);
  VGA_l076_g12526 : OAI22D0BWP7T port map(A1 => VGA_l076_n_66, A2 => VGA_l076_n_31, B1 => VGA_l076_n_47, B2 => VGA_x(2), ZN => VGA_l076_n_125);
  VGA_l076_g12527 : AN3D0BWP7T port map(A1 => VGA_l076_n_68, A2 => VGA_l076_n_75, A3 => VGA_l076_n_69, Z => VGA_l076_n_124);
  VGA_l076_g12528 : AN2D1BWP7T port map(A1 => VGA_l076_n_88, A2 => VGA_l076_n_68, Z => VGA_l076_n_123);
  VGA_l076_g12529 : AN2D1BWP7T port map(A1 => VGA_l076_n_89, A2 => VGA_l076_n_58, Z => VGA_l076_n_122);
  VGA_l076_g12530 : AOI221D0BWP7T port map(A1 => VGA_l076_n_61, A2 => VGA_draw_count10(0), B1 => VGA_l076_n_56, B2 => VGA_l076_n_25, C => VGA_l076_n_80, ZN => VGA_l076_n_112);
  VGA_l076_g12531 : AO222D0BWP7T port map(A1 => VGA_l076_n_61, A2 => VGA_l076_n_24, B1 => VGA_l076_n_55, B2 => VGA_l076_n_13, C1 => VGA_l076_n_53, C2 => VGA_l076_n_27, Z => VGA_l076_n_111);
  VGA_l076_g12532 : OAI22D0BWP7T port map(A1 => VGA_l076_n_45, A2 => VGA_l076_n_26, B1 => VGA_l076_n_46, B2 => VGA_l076_n_16, ZN => VGA_l076_n_110);
  VGA_l076_g12533 : MAOI22D0BWP7T port map(A1 => VGA_l076_n_50, A2 => VGA_l076_n_35, B1 => VGA_l076_n_50, B2 => VGA_l076_n_35, ZN => VGA_l076_n_109);
  VGA_l076_g12534 : OAI22D0BWP7T port map(A1 => VGA_l076_n_65, A2 => VGA_l076_n_15, B1 => VGA_l076_n_36, B2 => VGA_y(9), ZN => VGA_l076_n_108);
  VGA_l076_g12535 : AOI22D0BWP7T port map(A1 => VGA_l076_n_65, A2 => VGA_l076_n_15, B1 => VGA_l076_n_36, B2 => VGA_y(9), ZN => VGA_l076_n_107);
  VGA_l076_g12536 : MAOI22D0BWP7T port map(A1 => VGA_l076_n_48, A2 => VGA_l076_n_28, B1 => VGA_l076_n_48, B2 => VGA_l076_n_28, ZN => VGA_l076_n_106);
  VGA_l076_g12538 : MAOI22D0BWP7T port map(A1 => VGA_l076_n_38, A2 => VGA_l076_n_19, B1 => VGA_l076_n_38, B2 => VGA_l076_n_19, ZN => VGA_l076_n_116);
  VGA_l076_g12540 : MOAI22D0BWP7T port map(A1 => VGA_l076_n_38, A2 => VGA_l076_n_22, B1 => VGA_l076_n_38, B2 => VGA_l076_n_22, ZN => VGA_l076_n_115);
  VGA_l076_g12541 : MAOI22D0BWP7T port map(A1 => VGA_l076_n_37, A2 => VGA_l076_n_33, B1 => VGA_l076_n_37, B2 => VGA_l076_n_33, ZN => VGA_l076_n_114);
  VGA_l076_g12542 : MOAI22D0BWP7T port map(A1 => VGA_l076_n_37, A2 => VGA_l076_n_23, B1 => VGA_l076_n_37, B2 => VGA_l076_n_23, ZN => VGA_l076_n_113);
  VGA_l076_g12543 : AOI21D0BWP7T port map(A1 => VGA_l076_n_56, A2 => VGA_l076_n_24, B => VGA_l076_n_63, ZN => VGA_l076_n_99);
  VGA_l076_g12544 : NR2D0BWP7T port map(A1 => VGA_l076_n_44, A2 => VGA_l076_n_34, ZN => VGA_l076_n_98);
  VGA_l076_g12545 : IND2D0BWP7T port map(A1 => VGA_l076_n_46, B1 => x_pos_e6(5), ZN => VGA_l076_n_97);
  VGA_l076_g12546 : ND2D0BWP7T port map(A1 => VGA_l076_n_46, A2 => VGA_l076_n_16, ZN => VGA_l076_n_105);
  VGA_l076_g12547 : NR2D0BWP7T port map(A1 => VGA_l076_n_66, A2 => VGA_l076_n_31, ZN => VGA_l076_n_96);
  VGA_l076_g12548 : NR2D0BWP7T port map(A1 => VGA_l076_n_71, A2 => VGA_l076_n_41, ZN => VGA_l076_n_104);
  VGA_l076_g12550 : NR2D0BWP7T port map(A1 => VGA_l076_n_79, A2 => VGA_l076_n_78, ZN => VGA_l076_n_103);
  VGA_l076_g12551 : NR2D0BWP7T port map(A1 => VGA_l076_n_71, A2 => VGA_l076_n_82, ZN => VGA_l076_n_102);
  VGA_l076_g12552 : ND2D0BWP7T port map(A1 => VGA_l076_n_82, A2 => VGA_y(1), ZN => VGA_l076_n_101);
  VGA_l076_g12553 : IND2D0BWP7T port map(A1 => VGA_y(1), B1 => VGA_l076_n_41, ZN => VGA_l076_n_100);
  VGA_l076_g12554 : CKND1BWP7T port map(I => VGA_l076_n_90, ZN => VGA_l076_n_91);
  VGA_l076_g12555 : AOI21D0BWP7T port map(A1 => VGA_l076_n_59, A2 => VGA_l076_n_25, B => VGA_l076_n_73, ZN => VGA_l076_n_86);
  VGA_l076_g12556 : OAI21D0BWP7T port map(A1 => VGA_l076_n_56, A2 => VGA_l076_n_53, B => VGA_l076_n_24, ZN => VGA_l076_n_85);
  VGA_l076_g12557 : AO21D0BWP7T port map(A1 => VGA_l076_n_60, A2 => VGA_l076_n_54, B => VGA_l076_n_62, Z => VGA_l076_n_84);
  VGA_l076_g12558 : IAO21D0BWP7T port map(A1 => VGA_l076_n_60, A2 => VGA_l076_n_13, B => VGA_l076_n_55, ZN => VGA_l076_n_94);
  VGA_l076_g12559 : OAI21D0BWP7T port map(A1 => VGA_l076_n_52, A2 => VGA_draw_count10(1), B => VGA_l076_n_70, ZN => VGA_l076_n_93);
  VGA_l076_g12560 : AOI22D0BWP7T port map(A1 => VGA_l076_n_51, A2 => VGA_x(0), B1 => VGA_x(1), B2 => VGA_l076_n_6, ZN => VGA_l076_n_83);
  VGA_l076_g12561 : OA22D0BWP7T port map(A1 => VGA_l076_n_64, A2 => VGA_l076_n_12, B1 => VGA_l076_n_25, B2 => VGA_l076_n_0, Z => VGA_l076_n_92);
  VGA_l076_g12562 : OAI21D0BWP7T port map(A1 => VGA_l076_n_57, A2 => VGA_l076_n_13, B => VGA_l076_n_69, ZN => VGA_l076_n_90);
  VGA_l076_g12563 : AOI22D0BWP7T port map(A1 => VGA_l076_n_56, A2 => VGA_l076_n_13, B1 => VGA_l076_n_59, B2 => VGA_l076_n_24, ZN => VGA_l076_n_89);
  VGA_l076_g12564 : IAO21D0BWP7T port map(A1 => VGA_l076_n_0, A2 => VGA_l076_n_24, B => VGA_l076_n_79, ZN => VGA_l076_n_88);
  VGA_l076_g12565 : MOAI22D0BWP7T port map(A1 => VGA_l076_n_43, A2 => VGA_y(0), B1 => VGA_l076_n_43, B2 => VGA_y(0), ZN => VGA_l076_n_87);
  VGA_l076_g12568 : INVD0BWP7T port map(I => VGA_l076_n_41, ZN => VGA_l076_n_82);
  VGA_l076_g12569 : CKND1BWP7T port map(I => VGA_l076_n_26, ZN => VGA_l076_n_81);
  VGA_l076_g12570 : NR2D0BWP7T port map(A1 => VGA_l076_n_54, A2 => VGA_draw_count10(1), ZN => VGA_l076_n_80);
  VGA_l076_g12571 : INR2D0BWP7T port map(A1 => VGA_l076_n_63, B1 => VGA_l076_n_25, ZN => VGA_l076_n_79);
  VGA_l076_g12572 : NR2D0BWP7T port map(A1 => VGA_l076_n_0, A2 => VGA_draw_count10(1), ZN => VGA_l076_n_78);
  VGA_l076_g12573 : NR2D0BWP7T port map(A1 => VGA_l076_n_57, A2 => VGA_l076_n_29, ZN => VGA_l076_n_77);
  VGA_l076_g12574 : ND2D0BWP7T port map(A1 => VGA_l076_n_55, A2 => VGA_draw_count10(1), ZN => VGA_l076_n_76);
  VGA_l076_g12575 : ND2D0BWP7T port map(A1 => VGA_l076_n_53, A2 => VGA_l076_n_13, ZN => VGA_l076_n_75);
  VGA_l076_g12576 : ND2D0BWP7T port map(A1 => VGA_l076_n_53, A2 => VGA_draw_count10(1), ZN => VGA_l076_n_74);
  VGA_l076_g12577 : NR2D0BWP7T port map(A1 => VGA_l076_n_56, A2 => VGA_l076_n_59, ZN => VGA_l076_n_67);
  VGA_l076_g12578 : AN2D1BWP7T port map(A1 => VGA_l076_n_63, A2 => VGA_l076_n_27, Z => VGA_l076_n_73);
  VGA_l076_g12579 : NR2D0BWP7T port map(A1 => VGA_l076_n_52, A2 => VGA_l076_n_13, ZN => VGA_l076_n_72);
  VGA_l076_g12580 : ND2D0BWP7T port map(A1 => VGA_l076_n_40, A2 => VGA_l076_n_43, ZN => VGA_l076_n_71);
  VGA_l076_g12581 : IND2D0BWP7T port map(A1 => VGA_l076_n_62, B1 => VGA_l076_n_56, ZN => VGA_l076_n_70);
  VGA_l076_g12582 : ND2D0BWP7T port map(A1 => VGA_l076_n_63, A2 => VGA_l076_n_13, ZN => VGA_l076_n_69);
  VGA_l076_g12583 : IND2D0BWP7T port map(A1 => VGA_l076_n_62, B1 => VGA_l076_n_63, ZN => VGA_l076_n_68);
  VGA_l076_g12584 : INVD0BWP7T port map(I => VGA_l076_n_61, ZN => VGA_l076_n_60);
  VGA_l076_g12585 : INVD0BWP7T port map(I => VGA_l076_n_59, ZN => VGA_l076_n_58);
  VGA_l076_g12586 : INVD1BWP7T port map(I => VGA_l076_n_57, ZN => VGA_l076_n_56);
  VGA_l076_g12587 : INVD0BWP7T port map(I => VGA_l076_n_55, ZN => VGA_l076_n_54);
  VGA_l076_g12588 : INVD0BWP7T port map(I => VGA_l076_n_53, ZN => VGA_l076_n_52);
  VGA_l076_g12589 : IAO21D0BWP7T port map(A1 => VGA_x(1), A2 => VGA_l076_n_6, B => x_pos_e6(0), ZN => VGA_l076_n_51);
  VGA_l076_g12590 : OAI21D0BWP7T port map(A1 => VGA_l076_n_7, A2 => x_pos_e6(4), B => VGA_l076_n_26, ZN => VGA_l076_n_66);
  VGA_l076_g12591 : AOI21D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l076_n_5, B => VGA_l076_n_28, ZN => VGA_l076_n_65);
  VGA_l076_g12592 : IND2D0BWP7T port map(A1 => VGA_l076_n_30, B1 => VGA_draw_count10(4), ZN => VGA_l076_n_64);
  VGA_l076_g12593 : INR2D0BWP7T port map(A1 => VGA_draw_count10(4), B1 => VGA_l076_n_17, ZN => VGA_l076_n_63);
  VGA_l076_g12594 : INR2D0BWP7T port map(A1 => VGA_l076_n_29, B1 => VGA_l076_n_27, ZN => VGA_l076_n_62);
  VGA_l076_g12596 : NR2D0BWP7T port map(A1 => VGA_l076_n_14, A2 => VGA_draw_count10(4), ZN => VGA_l076_n_61);
  VGA_l076_g12597 : NR2D0BWP7T port map(A1 => VGA_l076_n_30, A2 => VGA_draw_count10(4), ZN => VGA_l076_n_59);
  VGA_l076_g12598 : IND2D0BWP7T port map(A1 => VGA_l076_n_14, B1 => VGA_draw_count10(4), ZN => VGA_l076_n_57);
  VGA_l076_g12599 : NR2D0BWP7T port map(A1 => VGA_l076_n_17, A2 => VGA_draw_count10(4), ZN => VGA_l076_n_55);
  VGA_l076_g12600 : NR2D0BWP7T port map(A1 => VGA_l076_n_18, A2 => VGA_draw_count10(4), ZN => VGA_l076_n_53);
  VGA_l076_g12601 : CKND1BWP7T port map(I => VGA_l076_n_43, ZN => VGA_l076_n_42);
  VGA_l076_g12602 : CKND1BWP7T port map(I => VGA_l076_n_40, ZN => VGA_l076_n_39);
  VGA_l076_g12603 : MOAI22D0BWP7T port map(A1 => VGA_y(8), A2 => y_pos_e6(8), B1 => VGA_y(8), B2 => y_pos_e6(8), ZN => VGA_l076_n_50);
  VGA_l076_g12604 : MOAI22D0BWP7T port map(A1 => VGA_x(7), A2 => x_pos_e6(7), B1 => VGA_x(7), B2 => x_pos_e6(7), ZN => VGA_l076_n_49);
  VGA_l076_g12605 : MOAI22D0BWP7T port map(A1 => VGA_y(7), A2 => y_pos_e6(7), B1 => VGA_y(7), B2 => y_pos_e6(7), ZN => VGA_l076_n_48);
  VGA_l076_g12606 : MAOI22D0BWP7T port map(A1 => VGA_x(3), A2 => x_pos_e6(3), B1 => VGA_x(3), B2 => x_pos_e6(3), ZN => VGA_l076_n_47);
  VGA_l076_g12607 : MOAI22D0BWP7T port map(A1 => VGA_x(6), A2 => x_pos_e6(6), B1 => VGA_x(6), B2 => x_pos_e6(6), ZN => VGA_l076_n_46);
  VGA_l076_g12608 : MOAI22D0BWP7T port map(A1 => VGA_x(5), A2 => x_pos_e6(5), B1 => VGA_x(5), B2 => x_pos_e6(5), ZN => VGA_l076_n_45);
  VGA_l076_g12609 : MAOI22D0BWP7T port map(A1 => VGA_y(5), A2 => y_pos_e6(5), B1 => VGA_y(5), B2 => y_pos_e6(5), ZN => VGA_l076_n_44);
  VGA_l076_g12610 : MOAI22D0BWP7T port map(A1 => VGA_y(1), A2 => y_pos_e6(1), B1 => VGA_y(1), B2 => y_pos_e6(1), ZN => VGA_l076_n_43);
  VGA_l076_g12611 : MOAI22D0BWP7T port map(A1 => VGA_y(2), A2 => y_pos_e6(2), B1 => VGA_y(2), B2 => y_pos_e6(2), ZN => VGA_l076_n_41);
  VGA_l076_g12612 : MOAI22D0BWP7T port map(A1 => VGA_y(0), A2 => y_pos_e6(0), B1 => VGA_y(0), B2 => y_pos_e6(0), ZN => VGA_l076_n_40);
  VGA_l076_g12613 : MAOI22D0BWP7T port map(A1 => VGA_y(4), A2 => y_pos_e6(4), B1 => VGA_y(4), B2 => y_pos_e6(4), ZN => VGA_l076_n_38);
  VGA_l076_g12614 : MOAI22D0BWP7T port map(A1 => VGA_y(3), A2 => y_pos_e6(3), B1 => VGA_y(3), B2 => y_pos_e6(3), ZN => VGA_l076_n_37);
  VGA_l076_g12615 : INVD1BWP7T port map(I => VGA_l076_n_25, ZN => VGA_l076_n_24);
  VGA_l076_g12616 : IND2D0BWP7T port map(A1 => VGA_y(8), B1 => y_pos_e6(8), ZN => VGA_l076_n_36);
  VGA_l076_g12617 : INR2D0BWP7T port map(A1 => y_pos_e6(7), B1 => VGA_y(7), ZN => VGA_l076_n_35);
  VGA_l076_g12618 : IND2D0BWP7T port map(A1 => y_pos_e6(4), B1 => VGA_y(4), ZN => VGA_l076_n_34);
  VGA_l076_g12619 : IND2D0BWP7T port map(A1 => y_pos_e6(2), B1 => VGA_y(2), ZN => VGA_l076_n_33);
  VGA_l076_g12620 : IND2D0BWP7T port map(A1 => x_pos_e6(6), B1 => VGA_x(6), ZN => VGA_l076_n_32);
  VGA_l076_g12621 : IND2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_e6(3), ZN => VGA_l076_n_31);
  VGA_l076_g12622 : ND2D0BWP7T port map(A1 => VGA_draw_count10(2), A2 => VGA_draw_count10(3), ZN => VGA_l076_n_30);
  VGA_l076_g12623 : ND2D0BWP7T port map(A1 => VGA_l076_n_3, A2 => VGA_draw_count10(0), ZN => VGA_l076_n_29);
  VGA_l076_g12624 : NR2D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_l076_n_5, ZN => VGA_l076_n_28);
  VGA_l076_g12625 : NR2D0BWP7T port map(A1 => VGA_l076_n_3, A2 => VGA_draw_count10(0), ZN => VGA_l076_n_27);
  VGA_l076_g12626 : ND2D0BWP7T port map(A1 => VGA_l076_n_7, A2 => x_pos_e6(4), ZN => VGA_l076_n_26);
  VGA_l076_g12627 : ND2D0BWP7T port map(A1 => VGA_draw_count10(1), A2 => VGA_draw_count10(0), ZN => VGA_l076_n_25);
  VGA_l076_g12629 : CKND1BWP7T port map(I => VGA_l076_n_13, ZN => VGA_l076_n_12);
  VGA_l076_g12630 : IND2D0BWP7T port map(A1 => VGA_y(4), B1 => y_pos_e6(4), ZN => VGA_l076_n_11);
  VGA_l076_g12631 : ND2D0BWP7T port map(A1 => VGA_l076_n_8, A2 => y_pos_e6(2), ZN => VGA_l076_n_23);
  VGA_l076_g12632 : NR2D0BWP7T port map(A1 => VGA_l076_n_9, A2 => y_pos_e6(3), ZN => VGA_l076_n_22);
  VGA_l076_g12633 : INR2D0BWP7T port map(A1 => x_pos_e6(7), B1 => VGA_x(7), ZN => VGA_l076_n_21);
  VGA_l076_g12634 : ND2D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_l076_n_10, ZN => VGA_l076_n_20);
  VGA_l076_g12635 : INR2D0BWP7T port map(A1 => y_pos_e6(3), B1 => VGA_y(3), ZN => VGA_l076_n_19);
  VGA_l076_g12636 : IND2D0BWP7T port map(A1 => VGA_draw_count10(2), B1 => VGA_draw_count10(3), ZN => VGA_l076_n_18);
  VGA_l076_g12637 : IND2D0BWP7T port map(A1 => VGA_draw_count10(3), B1 => VGA_draw_count10(2), ZN => VGA_l076_n_17);
  VGA_l076_g12638 : INR2D0BWP7T port map(A1 => VGA_x(5), B1 => x_pos_e6(5), ZN => VGA_l076_n_16);
  VGA_l076_g12639 : IND2D0BWP7T port map(A1 => y_pos_e6(5), B1 => VGA_y(5), ZN => VGA_l076_n_15);
  VGA_l076_g12640 : OR2D0BWP7T port map(A1 => VGA_draw_count10(2), A2 => VGA_draw_count10(3), Z => VGA_l076_n_14);
  VGA_l076_g12641 : NR2D0BWP7T port map(A1 => VGA_draw_count10(1), A2 => VGA_draw_count10(0), ZN => VGA_l076_n_13);
  VGA_l076_g12642 : CKND1BWP7T port map(I => x_pos_e6(8), ZN => VGA_l076_n_10);
  VGA_l076_g12643 : CKND1BWP7T port map(I => VGA_y(3), ZN => VGA_l076_n_9);
  VGA_l076_g12644 : CKND1BWP7T port map(I => VGA_y(2), ZN => VGA_l076_n_8);
  VGA_l076_g12645 : CKND1BWP7T port map(I => VGA_x(4), ZN => VGA_l076_n_7);
  VGA_l076_g12646 : CKND1BWP7T port map(I => x_pos_e6(1), ZN => VGA_l076_n_6);
  VGA_l076_g12647 : CKND1BWP7T port map(I => y_pos_e6(6), ZN => VGA_l076_n_5);
  VGA_l076_g12648 : CKND1BWP7T port map(I => y_pos_e6(1), ZN => VGA_l076_n_4);
  VGA_l076_g12649 : INVD0BWP7T port map(I => VGA_draw_count10(1), ZN => VGA_l076_n_3);
  VGA_l076_g2 : MUX2ND0BWP7T port map(I0 => VGA_y(3), I1 => VGA_l076_n_9, S => VGA_l076_n_38, ZN => VGA_l076_n_2);
  VGA_l076_g12650 : MUX2ND0BWP7T port map(I0 => VGA_l076_n_8, I1 => VGA_y(2), S => VGA_l076_n_37, ZN => VGA_l076_n_1);
  VGA_l076_g12651 : IND2D1BWP7T port map(A1 => VGA_l076_n_18, B1 => VGA_draw_count10(4), ZN => VGA_l076_n_0);
  VGA_l076_g12652 : INVD0BWP7T port map(I => VGA_l076_n_66, ZN => VGA_l076_n_95);
  VGA_l01_count_reg_8 : DFQD1BWP7T port map(CP => clk, D => VGA_l01_n_32, Q => VGA_x(8));
  VGA_l01_g630 : AO211D0BWP7T port map(A1 => VGA_l01_n_24, A2 => VGA_x(8), B => VGA_l01_n_29, C => reset, Z => VGA_l01_n_32);
  VGA_l01_g631 : AO211D0BWP7T port map(A1 => VGA_l01_n_19, A2 => VGA_x(7), B => VGA_l01_n_28, C => reset, Z => VGA_l01_n_31);
  VGA_l01_g633 : AO211D0BWP7T port map(A1 => VGA_l01_n_22, A2 => VGA_x(6), B => VGA_l01_n_27, C => reset, Z => VGA_l01_n_30);
  VGA_l01_g634 : NR4D0BWP7T port map(A1 => VGA_l01_n_22, A2 => VGA_l01_n_3, A3 => VGA_l01_n_5, A4 => VGA_x(8), ZN => VGA_l01_n_29);
  VGA_l01_g635 : OAI32D0BWP7T port map(A1 => VGA_x(7), A2 => VGA_l01_n_3, A3 => VGA_l01_n_22, B1 => VGA_l01_n_6, B2 => VGA_l01_n_7, ZN => VGA_l01_n_28);
  VGA_l01_count_reg_5 : DFQD1BWP7T port map(CP => clk, D => VGA_l01_n_26, Q => VGA_x(5));
  VGA_l01_g638 : NR2D0BWP7T port map(A1 => VGA_l01_n_22, A2 => VGA_x(6), ZN => VGA_l01_n_27);
  VGA_l01_g639 : AO211D0BWP7T port map(A1 => VGA_l01_n_20, A2 => VGA_x(5), B => VGA_l01_n_23, C => reset, Z => VGA_l01_n_26);
  VGA_l01_g640 : AO211D0BWP7T port map(A1 => VGA_l01_n_17, A2 => VGA_x(4), B => VGA_l01_n_21, C => reset, Z => VGA_l01_n_25);
  VGA_l01_g641 : AO211D0BWP7T port map(A1 => VGA_l01_n_3, A2 => VGA_x(5), B => VGA_l01_n_19, C => VGA_l01_n_5, Z => VGA_l01_n_24);
  VGA_l01_g642 : NR2D0BWP7T port map(A1 => VGA_l01_n_20, A2 => VGA_x(5), ZN => VGA_l01_n_23);
  VGA_l01_count_reg_3 : DFQD1BWP7T port map(CP => clk, D => VGA_l01_n_18, Q => VGA_x(3));
  VGA_l01_g644 : AOI211D0BWP7T port map(A1 => VGA_l01_n_8, A2 => VGA_l01_n_6, B => VGA_l01_n_17, C => VGA_x(4), ZN => VGA_l01_n_21);
  VGA_l01_g645 : IND2D0BWP7T port map(A1 => VGA_l01_n_20, B1 => VGA_x(5), ZN => VGA_l01_n_22);
  VGA_l01_g646 : IND2D0BWP7T port map(A1 => VGA_l01_n_17, B1 => VGA_x(4), ZN => VGA_l01_n_20);
  VGA_l01_g647 : AO211D0BWP7T port map(A1 => VGA_l01_n_14, A2 => VGA_x(3), B => VGA_l01_n_16, C => reset, Z => VGA_l01_n_18);
  VGA_l01_g648 : OR2D0BWP7T port map(A1 => VGA_l01_n_17, A2 => VGA_l01_n_11, Z => VGA_l01_n_19);
  VGA_l01_count_reg_2 : DFQD1BWP7T port map(CP => clk, D => VGA_l01_n_15, Q => VGA_x(2));
  VGA_l01_g650 : IND2D0BWP7T port map(A1 => VGA_l01_n_14, B1 => VGA_x(3), ZN => VGA_l01_n_17);
  VGA_l01_g651 : NR2D0BWP7T port map(A1 => VGA_l01_n_14, A2 => VGA_x(3), ZN => VGA_l01_n_16);
  VGA_l01_g652 : AO211D0BWP7T port map(A1 => VGA_l01_n_10, A2 => VGA_x(2), B => VGA_l01_n_13, C => reset, Z => VGA_l01_n_15);
  VGA_l01_count_reg_1 : DFQD1BWP7T port map(CP => clk, D => VGA_l01_n_12, Q => VGA_x(1));
  VGA_l01_g654 : IND2D0BWP7T port map(A1 => VGA_l01_n_10, B1 => VGA_x(2), ZN => VGA_l01_n_14);
  VGA_l01_g655 : NR2D0BWP7T port map(A1 => VGA_l01_n_10, A2 => VGA_x(2), ZN => VGA_l01_n_13);
  VGA_l01_g656 : AO211D0BWP7T port map(A1 => VGA_l01_n_2, A2 => VGA_x(1), B => VGA_l01_n_9, C => reset, Z => VGA_l01_n_12);
  VGA_l01_g657 : OAI222D0BWP7T port map(A1 => VGA_l01_n_4, A2 => VGA_x(6), B1 => VGA_x(5), B2 => VGA_l01_n_3, C1 => VGA_x(4), C2 => VGA_l01_n_3, ZN => VGA_l01_n_11);
  VGA_l01_count_reg_0 : DFKSND1BWP7T port map(CP => clk, D => reset, SN => VGA_x(0), Q => VGA_x(0), QN => VGA_l01_n_2);
  VGA_l01_g659 : NR2D0BWP7T port map(A1 => VGA_l01_n_2, A2 => VGA_x(1), ZN => VGA_l01_n_9);
  VGA_l01_g660 : ND2D0BWP7T port map(A1 => VGA_x(0), A2 => VGA_x(1), ZN => VGA_l01_n_10);
  VGA_l01_g661 : CKND1BWP7T port map(I => VGA_l01_n_7, ZN => VGA_l01_n_8);
  VGA_l01_g662 : ND2D0BWP7T port map(A1 => VGA_l01_n_3, A2 => VGA_x(7), ZN => VGA_l01_n_7);
  VGA_l01_g663 : INR2D0BWP7T port map(A1 => VGA_x(8), B1 => VGA_x(5), ZN => VGA_l01_n_6);
  VGA_l01_count_reg_7 : DFD1BWP7T port map(CP => clk, D => VGA_l01_n_31, Q => VGA_x(7), QN => VGA_l01_n_5);
  VGA_l01_count_reg_4 : DFD1BWP7T port map(CP => clk, D => VGA_l01_n_25, Q => VGA_x(4), QN => VGA_l01_n_4);
  VGA_l01_count_reg_6 : DFD1BWP7T port map(CP => clk, D => VGA_l01_n_30, Q => VGA_x(6), QN => VGA_l01_n_3);
  VGA_l02_count_reg_9 : DFQD1BWP7T port map(CP => clk, D => VGA_l02_n_40, Q => VGA_y(9));
  VGA_l02_g1038 : AO22D0BWP7T port map(A1 => VGA_l02_n_1, A2 => VGA_y(9), B1 => VGA_l02_n_23, B2 => VGA_l02_n_38, Z => VGA_l02_n_40);
  VGA_l02_g1039 : AO21D0BWP7T port map(A1 => VGA_l02_n_1, A2 => VGA_y(8), B => VGA_l02_n_37, Z => VGA_l02_n_39);
  VGA_l02_count_reg_7 : DFQD1BWP7T port map(CP => clk, D => VGA_l02_n_36, Q => VGA_y(7));
  VGA_l02_g1041 : OAI31D0BWP7T port map(A1 => VGA_y(9), A2 => VGA_l02_n_6, A3 => VGA_l02_n_32, B => VGA_l02_n_7, ZN => VGA_l02_n_38);
  VGA_l02_g1042 : NR3D0BWP7T port map(A1 => VGA_l02_n_32, A2 => VGA_l02_n_22, A3 => VGA_y(8), ZN => VGA_l02_n_37);
  VGA_l02_g1043 : MOAI22D0BWP7T port map(A1 => VGA_l02_n_33, A2 => VGA_l02_n_22, B1 => VGA_l02_n_15, B2 => VGA_y(7), ZN => VGA_l02_n_36);
  VGA_l02_g1047 : OAI22D0BWP7T port map(A1 => VGA_l02_n_30, A2 => VGA_l02_n_4, B1 => VGA_l02_n_22, B2 => VGA_l02_n_31, ZN => VGA_l02_n_35);
  VGA_l02_g1048 : OAI32D0BWP7T port map(A1 => VGA_y(5), A2 => VGA_l02_n_20, A3 => VGA_l02_n_22, B1 => VGA_l02_n_5, B2 => VGA_l02_n_30, ZN => VGA_l02_n_34);
  VGA_l02_g1049 : MAOI22D0BWP7T port map(A1 => VGA_l02_n_29, A2 => VGA_y(7), B1 => VGA_l02_n_29, B2 => VGA_y(7), ZN => VGA_l02_n_33);
  VGA_l02_count_reg_4 : DFQD1BWP7T port map(CP => clk, D => VGA_l02_n_28, Q => VGA_y(4));
  VGA_l02_g1051 : MAOI22D0BWP7T port map(A1 => VGA_l02_n_5, A2 => VGA_y(6), B1 => VGA_l02_n_27, B2 => VGA_y(6), ZN => VGA_l02_n_31);
  VGA_l02_g1052 : IND2D0BWP7T port map(A1 => VGA_l02_n_29, B1 => VGA_y(7), ZN => VGA_l02_n_32);
  VGA_l02_count_reg_1 : DFQD1BWP7T port map(CP => clk, D => VGA_l02_n_26, Q => VGA_y(1));
  VGA_l02_count_reg_3 : DFQD1BWP7T port map(CP => clk, D => VGA_l02_n_24, Q => VGA_y(3));
  VGA_l02_count_reg_2 : DFQD1BWP7T port map(CP => clk, D => VGA_l02_n_25, Q => VGA_y(2));
  VGA_l02_g1056 : MOAI22D0BWP7T port map(A1 => VGA_l02_n_22, A2 => VGA_l02_n_21, B1 => VGA_l02_n_15, B2 => VGA_y(4), ZN => VGA_l02_n_28);
  VGA_l02_g1057 : AOI21D0BWP7T port map(A1 => VGA_l02_n_23, A2 => VGA_l02_n_20, B => VGA_l02_n_15, ZN => VGA_l02_n_30);
  VGA_l02_g1058 : IND2D0BWP7T port map(A1 => VGA_l02_n_27, B1 => VGA_y(6), ZN => VGA_l02_n_29);
  VGA_l02_count_reg_0 : DFXQD1BWP7T port map(CP => clk, DA => VGA_l02_n_15, DB => VGA_l02_n_23, SA => VGA_y(0), Q => VGA_y(0));
  VGA_l02_g1060 : MOAI22D0BWP7T port map(A1 => VGA_l02_n_22, A2 => VGA_l02_n_0, B1 => VGA_l02_n_15, B2 => VGA_y(1), ZN => VGA_l02_n_26);
  VGA_l02_g1061 : IND2D0BWP7T port map(A1 => VGA_l02_n_20, B1 => VGA_y(5), ZN => VGA_l02_n_27);
  VGA_l02_g1062 : MOAI22D0BWP7T port map(A1 => VGA_l02_n_22, A2 => VGA_l02_n_14, B1 => VGA_l02_n_15, B2 => VGA_y(2), ZN => VGA_l02_n_25);
  VGA_l02_g1063 : MOAI22D0BWP7T port map(A1 => VGA_l02_n_22, A2 => VGA_l02_n_18, B1 => VGA_l02_n_15, B2 => VGA_y(3), ZN => VGA_l02_n_24);
  VGA_l02_g1064 : INVD1BWP7T port map(I => VGA_l02_n_23, ZN => VGA_l02_n_22);
  VGA_l02_g1065 : NR3D0BWP7T port map(A1 => VGA_l02_n_19, A2 => VGA_l02_n_12, A3 => reset, ZN => VGA_l02_n_23);
  VGA_l02_g1066 : MAOI22D0BWP7T port map(A1 => VGA_l02_n_17, A2 => VGA_y(4), B1 => VGA_l02_n_17, B2 => VGA_y(4), ZN => VGA_l02_n_21);
  VGA_l02_g1067 : IND2D0BWP7T port map(A1 => VGA_l02_n_17, B1 => VGA_y(4), ZN => VGA_l02_n_20);
  VGA_l02_g1068 : NR4D0BWP7T port map(A1 => VGA_l02_n_16, A2 => VGA_y(6), A3 => VGA_y(7), A4 => VGA_y(5), ZN => VGA_l02_n_19);
  VGA_l02_g1069 : MAOI22D0BWP7T port map(A1 => VGA_l02_n_13, A2 => VGA_y(3), B1 => VGA_l02_n_13, B2 => VGA_y(3), ZN => VGA_l02_n_18);
  VGA_l02_g1070 : IND2D0BWP7T port map(A1 => VGA_l02_n_13, B1 => VGA_y(3), ZN => VGA_l02_n_17);
  VGA_l02_g1071 : IND4D0BWP7T port map(A1 => VGA_y(4), B1 => VGA_y(2), B2 => VGA_y(3), B3 => VGA_l02_n_11, ZN => VGA_l02_n_16);
  VGA_l02_g1073 : INR2D0BWP7T port map(A1 => VGA_l02_n_12, B1 => reset, ZN => VGA_l02_n_15);
  VGA_l02_g1074 : MAOI22D0BWP7T port map(A1 => VGA_l02_n_8, A2 => VGA_y(2), B1 => VGA_l02_n_8, B2 => VGA_y(2), ZN => VGA_l02_n_14);
  VGA_l02_g1075 : IND2D0BWP7T port map(A1 => VGA_l02_n_8, B1 => VGA_y(2), ZN => VGA_l02_n_13);
  VGA_l02_g1076 : IND4D0BWP7T port map(A1 => VGA_l02_n_10, B1 => VGA_x(1), B2 => VGA_x(2), B3 => VGA_l02_n_9, ZN => VGA_l02_n_12);
  VGA_l02_g1077 : NR3D0BWP7T port map(A1 => VGA_l02_n_7, A2 => VGA_y(0), A3 => VGA_y(1), ZN => VGA_l02_n_11);
  VGA_l02_g1078 : ND3D0BWP7T port map(A1 => VGA_x(8), A2 => VGA_x(7), A3 => VGA_x(0), ZN => VGA_l02_n_10);
  VGA_l02_g1079 : INR4D0BWP7T port map(A1 => VGA_x(3), B1 => VGA_x(6), B2 => VGA_x(4), B3 => VGA_x(5), ZN => VGA_l02_n_9);
  VGA_l02_g1081 : ND2D0BWP7T port map(A1 => VGA_y(0), A2 => VGA_y(1), ZN => VGA_l02_n_8);
  VGA_l02_g1082 : ND2D0BWP7T port map(A1 => VGA_l02_n_6, A2 => VGA_y(9), ZN => VGA_l02_n_7);
  VGA_l02_g2 : AO21D0BWP7T port map(A1 => VGA_l02_n_32, A2 => VGA_l02_n_23, B => VGA_l02_n_15, Z => VGA_l02_n_1);
  VGA_l02_g1092 : XNR2D1BWP7T port map(A1 => VGA_y(1), A2 => VGA_y(0), ZN => VGA_l02_n_0);
  VGA_l02_count_reg_8 : DFD1BWP7T port map(CP => clk, D => VGA_l02_n_39, Q => VGA_y(8), QN => VGA_l02_n_6);
  VGA_l02_count_reg_5 : DFD1BWP7T port map(CP => clk, D => VGA_l02_n_34, Q => VGA_y(5), QN => VGA_l02_n_5);
  VGA_l02_count_reg_6 : DFD1BWP7T port map(CP => clk, D => VGA_l02_n_35, Q => VGA_y(6), QN => VGA_l02_n_4);
  VGA_l03_hold_reg : DFD1BWP7T port map(CP => clk, D => VGA_l03_n_11, Q => UNCONNECTED, QN => VGA_l03_n_13);
  VGA_l03_g308 : INVD4BWP7T port map(I => VGA_l03_n_13, ZN => h_sync);
  VGA_l03_vold_reg : DFD1BWP7T port map(CP => clk, D => VGA_l03_n_35, Q => UNCONNECTED0, QN => VGA_l03_n_12);
  VGA_l03_g310 : INVD4BWP7T port map(I => VGA_l03_n_12, ZN => v_sync);
  VGA_l03_g311 : NR2D0BWP7T port map(A1 => VGA_l03_n_36, A2 => reset, ZN => VGA_l03_n_11);
  VGA_l03_g314 : IIND4D0BWP7T port map(A1 => VGA_y(6), A2 => VGA_y(2), B1 => VGA_l03_n_3, B2 => VGA_l03_n_6, ZN => VGA_l03_n_8);
  VGA_l03_g315 : OAI21D0BWP7T port map(A1 => VGA_l03_n_4, A2 => VGA_x(8), B => VGA_l03_n_2, ZN => VGA_l03_n_7);
  VGA_l03_g316 : NR3D0BWP7T port map(A1 => VGA_y(3), A2 => VGA_y(9), A3 => VGA_y(1), ZN => VGA_l03_n_6);
  VGA_l03_g317 : NR3D0BWP7T port map(A1 => VGA_x(6), A2 => VGA_x(4), A3 => VGA_x(5), ZN => VGA_l03_n_5);
  VGA_l03_g318 : AOI21D0BWP7T port map(A1 => VGA_x(4), A2 => VGA_x(5), B => VGA_x(6), ZN => VGA_l03_n_4);
  VGA_l03_g319 : NR4D0BWP7T port map(A1 => VGA_y(7), A2 => VGA_y(8), A3 => VGA_y(5), A4 => VGA_y(4), ZN => VGA_l03_n_3);
  VGA_l03_g320 : XNR2D1BWP7T port map(A1 => VGA_x(8), A2 => VGA_x(7), ZN => VGA_l03_n_2);
  VGA_l03_g2 : INR2D1BWP7T port map(A1 => VGA_l03_n_8, B1 => reset, ZN => VGA_l03_n_35);
  VGA_l03_g325 : AOI21D0BWP7T port map(A1 => VGA_l03_n_5, A2 => VGA_x(8), B => VGA_l03_n_7, ZN => VGA_l03_n_36);
  Enemy_spawning_en11_decider_reg : DFQD1BWP7T port map(CP => clk, D => Enemy_spawning_en11_n_3, Q => spawn_or_not_e1);
  Enemy_spawning_en11_g143 : NR4D0BWP7T port map(A1 => Enemy_spawning_en11_n_2, A2 => Enemy_spawning_en11_n_1, A3 => Enemy_spawning_en11_n_0, A4 => e_1, ZN => Enemy_spawning_en11_n_3);
  Enemy_spawning_en11_g144 : ND4D0BWP7T port map(A1 => y_e_spawn_3(7), A2 => y_e_spawn_4(7), A3 => y_e_spawn_2(3), A4 => y_e_spawn_2(1), ZN => Enemy_spawning_en11_n_2);
  Enemy_spawning_en11_g145 : ND2D0BWP7T port map(A1 => y_e_spawn_5(8), A2 => y_e_spawn_2(7), ZN => Enemy_spawning_en11_n_1);
  Enemy_spawning_en11_g146 : ND2D0BWP7T port map(A1 => y_e_spawn_3(3), A2 => n_5, ZN => Enemy_spawning_en11_n_0);
  Enemy_spawning_en21_decider_reg : DFQD1BWP7T port map(CP => clk, D => Enemy_spawning_en21_n_3, Q => spawn_or_not_e2);
  Enemy_spawning_en21_g143 : NR4D0BWP7T port map(A1 => Enemy_spawning_en21_n_2, A2 => Enemy_spawning_en21_n_1, A3 => Enemy_spawning_en21_n_0, A4 => e_2, ZN => Enemy_spawning_en21_n_3);
  Enemy_spawning_en21_g144 : ND4D0BWP7T port map(A1 => y_e_spawn_1(4), A2 => y_e_spawn_1(5), A3 => y_e_spawn_2(1), A4 => y_e_spawn_1(2), ZN => Enemy_spawning_en21_n_2);
  Enemy_spawning_en21_g145 : ND2D0BWP7T port map(A1 => y_e_spawn_1(8), A2 => y_e_spawn_2(7), ZN => Enemy_spawning_en21_n_1);
  Enemy_spawning_en21_g146 : ND2D0BWP7T port map(A1 => y_e_spawn_1(1), A2 => n_5, ZN => Enemy_spawning_en21_n_0);
  Enemy_spawning_en31_decider_reg : DFQD1BWP7T port map(CP => clk, D => Enemy_spawning_en31_n_3, Q => spawn_or_not_e3);
  Enemy_spawning_en31_g143 : NR4D0BWP7T port map(A1 => Enemy_spawning_en31_n_2, A2 => Enemy_spawning_en31_n_1, A3 => Enemy_spawning_en31_n_0, A4 => e_3, ZN => Enemy_spawning_en31_n_3);
  Enemy_spawning_en31_g144 : ND4D0BWP7T port map(A1 => y_e_spawn_1(3), A2 => y_e_spawn_1(5), A3 => y_e_spawn_2(1), A4 => y_e_spawn_1(2), ZN => Enemy_spawning_en31_n_2);
  Enemy_spawning_en31_g145 : ND2D0BWP7T port map(A1 => y_e_spawn_5(8), A2 => y_e_spawn_1(8), ZN => Enemy_spawning_en31_n_1);
  Enemy_spawning_en31_g146 : ND2D0BWP7T port map(A1 => y_e_spawn_1(0), A2 => n_5, ZN => Enemy_spawning_en31_n_0);
  Enemy_spawning_en41_decider_reg : DFQD1BWP7T port map(CP => clk, D => Enemy_spawning_en41_n_3, Q => spawn_or_not_e4);
  Enemy_spawning_en41_g143 : NR4D0BWP7T port map(A1 => Enemy_spawning_en41_n_2, A2 => Enemy_spawning_en41_n_1, A3 => Enemy_spawning_en41_n_0, A4 => e_4, ZN => Enemy_spawning_en41_n_3);
  Enemy_spawning_en41_g144 : ND4D0BWP7T port map(A1 => y_e_spawn_1(4), A2 => y_e_spawn_3(7), A3 => y_e_spawn_1(8), A4 => y_e_spawn_1(3), ZN => Enemy_spawning_en41_n_2);
  Enemy_spawning_en41_g145 : ND2D0BWP7T port map(A1 => y_e_spawn_1(7), A2 => y_e_spawn_4(7), ZN => Enemy_spawning_en41_n_1);
  Enemy_spawning_en41_g146 : ND2D0BWP7T port map(A1 => y_e_spawn_1(0), A2 => n_5, ZN => Enemy_spawning_en41_n_0);
  VGA_l041_count_reg_2 : DFCNQD1BWP7T port map(CDN => VGA_l041_n_0, CP => clk, D => VGA_l041_n_6, Q => VGA_draw_count1(2));
  VGA_l041_g59 : INR2D0BWP7T port map(A1 => VGA_enable1, B1 => VGA_l041_n_5, ZN => VGA_l041_n_6);
  VGA_l041_count_reg_1 : DFCNQD1BWP7T port map(CDN => VGA_l041_n_0, CP => clk, D => VGA_l041_n_4, Q => VGA_draw_count1(1));
  VGA_l041_g61 : MAOI22D0BWP7T port map(A1 => VGA_l041_n_1, A2 => VGA_draw_count1(2), B1 => VGA_l041_n_1, B2 => VGA_draw_count1(2), ZN => VGA_l041_n_5);
  VGA_l041_g62 : INR2D0BWP7T port map(A1 => VGA_enable1, B1 => VGA_l041_n_3, ZN => VGA_l041_n_4);
  VGA_l041_count_reg_0 : DFCNQD1BWP7T port map(CDN => VGA_l041_n_0, CP => clk, D => VGA_l041_n_2, Q => VGA_draw_count1(0));
  VGA_l041_g64 : XNR2D1BWP7T port map(A1 => VGA_draw_count1(0), A2 => VGA_draw_count1(1), ZN => VGA_l041_n_3);
  VGA_l041_g65 : INR2D0BWP7T port map(A1 => VGA_enable1, B1 => VGA_draw_count1(0), ZN => VGA_l041_n_2);
  VGA_l041_g66 : ND2D0BWP7T port map(A1 => VGA_draw_count1(0), A2 => VGA_draw_count1(1), ZN => VGA_l041_n_1);
  VGA_l041_g67 : INVD0BWP7T port map(I => reset, ZN => VGA_l041_n_0);
  VGA_l06_g13497 : IND4D0BWP7T port map(A1 => VGA_l06_n_286, B1 => VGA_l06_n_298, B2 => VGA_l06_n_295, B3 => VGA_l06_n_323, ZN => VGA_b4);
  VGA_l06_g13498 : ND3D0BWP7T port map(A1 => VGA_l06_n_322, A2 => VGA_l06_n_293, A3 => VGA_l06_n_281, ZN => VGA_g4);
  VGA_l06_g13499 : NR4D0BWP7T port map(A1 => VGA_l06_n_319, A2 => VGA_l06_n_267, A3 => VGA_l06_n_253, A4 => VGA_l06_n_280, ZN => VGA_l06_n_323);
  VGA_l06_g13500 : AOI211D0BWP7T port map(A1 => VGA_l06_n_240, A2 => VGA_l06_n_135, B => VGA_l06_n_320, C => VGA_l06_n_297, ZN => VGA_l06_n_322);
  VGA_l06_g13501 : IND4D0BWP7T port map(A1 => VGA_l06_n_318, B1 => VGA_l06_n_265, B2 => VGA_l06_n_255, B3 => VGA_l06_n_275, ZN => VGA_r4);
  VGA_l06_g13502 : ND4D0BWP7T port map(A1 => VGA_l06_n_314, A2 => VGA_l06_n_306, A3 => VGA_l06_n_303, A4 => VGA_l06_n_282, ZN => VGA_l06_n_320);
  VGA_l06_g13503 : IND4D0BWP7T port map(A1 => VGA_l06_n_296, B1 => VGA_l06_n_258, B2 => VGA_l06_n_294, B3 => VGA_l06_n_316, ZN => VGA_l06_n_319);
  VGA_l06_g13504 : OAI211D0BWP7T port map(A1 => VGA_l06_n_217, A2 => VGA_l06_n_302, B => VGA_l06_n_315, C => VGA_l06_n_306, ZN => VGA_l06_n_318);
  VGA_l06_g13505 : IND3D0BWP7T port map(A1 => VGA_l06_n_240, B1 => VGA_l06_n_261, B2 => VGA_l06_n_312, ZN => VGA_enable4);
  VGA_l06_g13506 : NR4D0BWP7T port map(A1 => VGA_l06_n_313, A2 => VGA_l06_n_284, A3 => VGA_l06_n_239, A4 => VGA_l06_n_233, ZN => VGA_l06_n_316);
  VGA_l06_g13507 : IINR4D0BWP7T port map(A1 => VGA_l06_n_303, A2 => VGA_l06_n_282, B1 => VGA_l06_n_308, B2 => VGA_l06_n_301, ZN => VGA_l06_n_315);
  VGA_l06_g13508 : AOI211D0BWP7T port map(A1 => VGA_l06_n_271, A2 => VGA_l06_n_176, B => VGA_l06_n_311, C => VGA_l06_n_288, ZN => VGA_l06_n_314);
  VGA_l06_g13509 : OAI211D0BWP7T port map(A1 => VGA_l06_n_193, A2 => VGA_l06_n_260, B => VGA_l06_n_310, C => VGA_l06_n_266, ZN => VGA_l06_n_313);
  VGA_l06_g13510 : AOI211D0BWP7T port map(A1 => VGA_l06_n_307, A2 => VGA_l06_n_216, B => VGA_l06_n_232, C => VGA_l06_n_241, ZN => VGA_l06_n_312);
  VGA_l06_g13511 : ND4D0BWP7T port map(A1 => VGA_l06_n_309, A2 => VGA_l06_n_289, A3 => VGA_l06_n_254, A4 => VGA_l06_n_251, ZN => VGA_l06_n_311);
  VGA_l06_g13512 : NR4D0BWP7T port map(A1 => VGA_l06_n_305, A2 => VGA_l06_n_291, A3 => VGA_l06_n_230, A4 => VGA_l06_n_257, ZN => VGA_l06_n_310);
  VGA_l06_g13513 : AOI211D0BWP7T port map(A1 => VGA_l06_n_269, A2 => VGA_l06_n_195, B => VGA_l06_n_300, C => VGA_l06_n_299, ZN => VGA_l06_n_309);
  VGA_l06_g13514 : OAI211D0BWP7T port map(A1 => VGA_l06_n_120, A2 => VGA_l06_n_245, B => VGA_l06_n_304, C => VGA_l06_n_285, ZN => VGA_l06_n_308);
  VGA_l06_g13515 : IND4D0BWP7T port map(A1 => VGA_l06_n_268, B1 => VGA_l06_n_5, B2 => VGA_l06_n_235, B3 => VGA_l06_n_283, ZN => VGA_l06_n_307);
  VGA_l06_g13516 : OAI211D0BWP7T port map(A1 => VGA_l06_n_201, A2 => VGA_l06_n_263, B => VGA_l06_n_279, C => VGA_l06_n_256, ZN => VGA_l06_n_305);
  VGA_l06_g13517 : AOI221D0BWP7T port map(A1 => VGA_l06_n_269, A2 => VGA_l06_n_173, B1 => VGA_l06_n_270, B2 => VGA_l06_n_15, C => VGA_l06_n_299, ZN => VGA_l06_n_304);
  VGA_l06_g13518 : ND2D0BWP7T port map(A1 => VGA_l06_n_292, A2 => VGA_l06_n_13, ZN => VGA_l06_n_306);
  VGA_l06_g13519 : AOI22D0BWP7T port map(A1 => VGA_l06_n_290, A2 => VGA_l06_n_80, B1 => VGA_l06_n_268, B2 => VGA_l06_n_86, ZN => VGA_l06_n_302);
  VGA_l06_g13520 : ND4D0BWP7T port map(A1 => VGA_l06_n_274, A2 => VGA_l06_n_278, A3 => VGA_l06_n_252, A4 => VGA_l06_n_287, ZN => VGA_l06_n_301);
  VGA_l06_g13521 : OAI211D0BWP7T port map(A1 => VGA_l06_n_211, A2 => VGA_l06_n_6, B => VGA_l06_n_277, C => VGA_l06_n_264, ZN => VGA_l06_n_300);
  VGA_l06_g13522 : AOI22D0BWP7T port map(A1 => VGA_l06_n_276, A2 => VGA_l06_n_216, B1 => VGA_l06_n_271, B2 => VGA_l06_n_186, ZN => VGA_l06_n_303);
  VGA_l06_g13523 : AOI22D0BWP7T port map(A1 => VGA_l06_n_206, A2 => VGA_l06_n_271, B1 => VGA_l06_n_241, B2 => VGA_l06_n_115, ZN => VGA_l06_n_298);
  VGA_l06_g13524 : NR3D0BWP7T port map(A1 => VGA_l06_n_273, A2 => VGA_l06_n_217, A3 => VGA_l06_n_116, ZN => VGA_l06_n_297);
  VGA_l06_g13525 : OAI33D0BWP7T port map(A1 => VGA_l06_n_184, A2 => VGA_l06_n_217, A3 => VGA_l06_n_235, B1 => VGA_l06_n_164, B2 => VGA_l06_n_179, B3 => VGA_l06_n_228, ZN => VGA_l06_n_296);
  VGA_l06_g13526 : AO22D0BWP7T port map(A1 => VGA_l06_n_270, A2 => VGA_l06_n_166, B1 => VGA_l06_n_158, B2 => VGA_l06_n_269, Z => VGA_l06_n_299);
  VGA_l06_g13527 : MAOI22D0BWP7T port map(A1 => VGA_l06_n_240, A2 => VGA_l06_n_154, B1 => VGA_l06_n_273, B2 => VGA_l06_n_225, ZN => VGA_l06_n_295);
  VGA_l06_g13528 : MAOI22D0BWP7T port map(A1 => VGA_l06_n_248, A2 => VGA_l06_n_182, B1 => VGA_l06_n_261, B2 => VGA_l06_n_12, ZN => VGA_l06_n_294);
  VGA_l06_g13529 : AOI22D0BWP7T port map(A1 => VGA_l06_n_268, A2 => VGA_l06_n_226, B1 => VGA_l06_n_244, B2 => VGA_l06_n_154, ZN => VGA_l06_n_293);
  VGA_l06_g13530 : OAI22D0BWP7T port map(A1 => VGA_l06_n_261, A2 => VGA_l06_n_118, B1 => VGA_l06_n_249, B2 => VGA_l06_n_88, ZN => VGA_l06_n_292);
  VGA_l06_g13531 : OA21D0BWP7T port map(A1 => VGA_l06_n_202, A2 => VGA_l06_n_158, B => VGA_l06_n_269, Z => VGA_l06_n_291);
  VGA_l06_g13532 : IND2D0BWP7T port map(A1 => VGA_l06_n_268, B1 => VGA_l06_n_273, ZN => VGA_l06_n_290);
  VGA_l06_g13533 : IND2D0BWP7T port map(A1 => VGA_l06_n_263, B1 => VGA_l06_n_207, ZN => VGA_l06_n_289);
  VGA_l06_g13534 : AOI31D0BWP7T port map(A1 => VGA_l06_n_3, A2 => VGA_l06_n_129, A3 => VGA_l06_n_123, B => VGA_l06_n_260, ZN => VGA_l06_n_288);
  VGA_l06_g13535 : IOA21D0BWP7T port map(A1 => VGA_l06_n_180, A2 => VGA_l06_n_120, B => VGA_l06_n_271, ZN => VGA_l06_n_287);
  VGA_l06_g13536 : NR3D0BWP7T port map(A1 => VGA_l06_n_237, A2 => VGA_l06_n_217, A3 => VGA_l06_n_136, ZN => VGA_l06_n_286);
  VGA_l06_g13537 : OAI31D0BWP7T port map(A1 => VGA_l06_n_31, A2 => VGA_l06_n_84, A3 => VGA_l06_n_199, B => VGA_l06_n_272, ZN => VGA_l06_n_285);
  VGA_l06_g13538 : AOI21D0BWP7T port map(A1 => VGA_l06_n_193, A2 => VGA_l06_n_159, B => VGA_l06_n_6, ZN => VGA_l06_n_284);
  VGA_l06_g13539 : NR3D0BWP7T port map(A1 => VGA_l06_n_231, A2 => VGA_l06_n_236, A3 => VGA_l06_n_222, ZN => VGA_l06_n_283);
  VGA_l06_g13540 : AOI22D0BWP7T port map(A1 => VGA_l06_n_242, A2 => VGA_l06_n_190, B1 => VGA_l06_n_241, B2 => VGA_l06_n_91, ZN => VGA_l06_n_281);
  VGA_l06_g13541 : AOI211D0BWP7T port map(A1 => VGA_l06_n_136, A2 => VGA_l06_n_77, B => VGA_l06_n_238, C => VGA_l06_n_217, ZN => VGA_l06_n_280);
  VGA_l06_g13542 : OAI21D0BWP7T port map(A1 => VGA_l06_n_205, A2 => VGA_l06_n_192, B => VGA_l06_n_270, ZN => VGA_l06_n_279);
  VGA_l06_g13543 : OAI21D0BWP7T port map(A1 => VGA_l06_n_154, A2 => VGA_l06_n_147, B => VGA_l06_n_259, ZN => VGA_l06_n_278);
  VGA_l06_g13544 : OAI21D0BWP7T port map(A1 => VGA_l06_n_183, A2 => VGA_l06_n_128, B => VGA_l06_n_270, ZN => VGA_l06_n_277);
  VGA_l06_g13545 : OAI22D0BWP7T port map(A1 => VGA_l06_n_5, A2 => VGA_l06_n_78, B1 => VGA_l06_n_235, B2 => VGA_l06_n_126, ZN => VGA_l06_n_276);
  VGA_l06_g13546 : AOI22D0BWP7T port map(A1 => VGA_l06_n_244, A2 => VGA_l06_n_155, B1 => VGA_l06_n_240, B2 => VGA_l06_n_137, ZN => VGA_l06_n_275);
  VGA_l06_g13547 : OAI21D0BWP7T port map(A1 => VGA_l06_n_176, A2 => VGA_l06_n_173, B => VGA_l06_n_262, ZN => VGA_l06_n_274);
  VGA_l06_g13548 : MAOI22D0BWP7T port map(A1 => VGA_l06_n_250, A2 => VGA_l06_n_181, B1 => VGA_l06_n_228, B2 => VGA_l06_n_203, ZN => VGA_l06_n_282);
  VGA_l06_g13549 : INVD0BWP7T port map(I => VGA_l06_n_6, ZN => VGA_l06_n_272);
  VGA_l06_g13550 : INR2D0BWP7T port map(A1 => VGA_l06_n_244, B1 => VGA_l06_n_185, ZN => VGA_l06_n_267);
  VGA_l06_g13551 : OAI21D0BWP7T port map(A1 => VGA_l06_n_181, A2 => VGA_l06_n_143, B => VGA_l06_n_246, ZN => VGA_l06_n_266);
  VGA_l06_g13552 : OAI21D0BWP7T port map(A1 => VGA_l06_n_161, A2 => VGA_l06_n_165, B => VGA_l06_n_242, ZN => VGA_l06_n_265);
  VGA_l06_g13553 : OAI31D0BWP7T port map(A1 => VGA_l06_n_144, A2 => VGA_l06_n_183, A3 => VGA_l06_n_176, B => VGA_l06_n_234, ZN => VGA_l06_n_264);
  VGA_l06_g13554 : AOI21D0BWP7T port map(A1 => VGA_l06_n_219, A2 => VGA_l06_n_178, B => VGA_l06_n_236, ZN => VGA_l06_n_273);
  VGA_l06_g13556 : NR4D0BWP7T port map(A1 => VGA_l06_n_215, A2 => VGA_l06_n_217, A3 => VGA_l06_n_47, A4 => VGA_l06_n_59, ZN => VGA_l06_n_271);
  VGA_l06_g13557 : NR2D0BWP7T port map(A1 => VGA_l06_n_247, A2 => VGA_l06_n_156, ZN => VGA_l06_n_270);
  VGA_l06_g13558 : NR2D0BWP7T port map(A1 => VGA_l06_n_247, A2 => VGA_l06_n_149, ZN => VGA_l06_n_269);
  VGA_l06_g13559 : ND2D0BWP7T port map(A1 => VGA_l06_n_238, A2 => VGA_l06_n_237, ZN => VGA_l06_n_268);
  VGA_l06_g13560 : CKND1BWP7T port map(I => VGA_l06_n_262, ZN => VGA_l06_n_263);
  VGA_l06_g13561 : CKND1BWP7T port map(I => VGA_l06_n_259, ZN => VGA_l06_n_260);
  VGA_l06_g13562 : OAI21D0BWP7T port map(A1 => VGA_l06_n_190, A2 => VGA_l06_n_121, B => VGA_l06_n_242, ZN => VGA_l06_n_258);
  VGA_l06_g13563 : OA21D0BWP7T port map(A1 => VGA_l06_n_170, A2 => VGA_l06_n_87, B => VGA_l06_n_250, Z => VGA_l06_n_257);
  VGA_l06_g13564 : OAI31D0BWP7T port map(A1 => VGA_l06_n_110, A2 => VGA_l06_n_192, A3 => VGA_l06_n_194, B => VGA_l06_n_234, ZN => VGA_l06_n_256);
  VGA_l06_g13565 : OAI21D0BWP7T port map(A1 => VGA_l06_n_155, A2 => VGA_l06_n_79, B => VGA_l06_n_243, ZN => VGA_l06_n_255);
  VGA_l06_g13566 : OAI21D0BWP7T port map(A1 => VGA_l06_n_154, A2 => VGA_l06_n_79, B => VGA_l06_n_243, ZN => VGA_l06_n_254);
  VGA_l06_g13567 : OA21D0BWP7T port map(A1 => VGA_l06_n_190, A2 => VGA_l06_n_90, B => VGA_l06_n_243, Z => VGA_l06_n_253);
  VGA_l06_g13568 : OAI31D0BWP7T port map(A1 => VGA_l06_n_15, A2 => VGA_l06_n_130, A3 => VGA_l06_n_191, B => VGA_l06_n_234, ZN => VGA_l06_n_252);
  VGA_l06_g13569 : OAI21D0BWP7T port map(A1 => VGA_l06_n_181, A2 => VGA_l06_n_76, B => VGA_l06_n_246, ZN => VGA_l06_n_251);
  VGA_l06_g13570 : NR3D0BWP7T port map(A1 => VGA_l06_n_229, A2 => VGA_l06_n_163, A3 => VGA_l06_n_96, ZN => VGA_l06_n_262);
  VGA_l06_g13571 : OR3D0BWP7T port map(A1 => VGA_l06_n_98, A2 => VGA_l06_n_149, A3 => VGA_l06_n_228, Z => VGA_l06_n_261);
  VGA_l06_g13572 : NR3D0BWP7T port map(A1 => VGA_l06_n_229, A2 => VGA_l06_n_1, A3 => VGA_l06_n_96, ZN => VGA_l06_n_259);
  VGA_l06_g13573 : CKND1BWP7T port map(I => VGA_l06_n_248, ZN => VGA_l06_n_249);
  VGA_l06_g13575 : INVD0BWP7T port map(I => VGA_l06_n_246, ZN => VGA_l06_n_245);
  VGA_l06_g13576 : AOI211D0BWP7T port map(A1 => VGA_l06_n_168, A2 => VGA_l06_n_169, B => VGA_l06_n_228, C => VGA_l06_n_140, ZN => VGA_l06_n_239);
  VGA_l06_g13577 : NR4D0BWP7T port map(A1 => VGA_l06_n_217, A2 => VGA_l06_n_213, A3 => VGA_l06_n_134, A4 => VGA_l06_n_60, ZN => VGA_l06_n_250);
  VGA_l06_g13578 : NR2D0BWP7T port map(A1 => VGA_l06_n_228, A2 => VGA_l06_n_139, ZN => VGA_l06_n_248);
  VGA_l06_g13579 : IND2D0BWP7T port map(A1 => VGA_l06_n_229, B1 => VGA_l06_n_98, ZN => VGA_l06_n_247);
  VGA_l06_g13580 : NR2D0BWP7T port map(A1 => VGA_l06_n_229, A2 => VGA_l06_n_174, ZN => VGA_l06_n_246);
  VGA_l06_g13581 : NR2D0BWP7T port map(A1 => VGA_l06_n_224, A2 => VGA_l06_n_179, ZN => VGA_l06_n_244);
  VGA_l06_g13582 : NR2D0BWP7T port map(A1 => VGA_l06_n_224, A2 => VGA_l06_n_169, ZN => VGA_l06_n_243);
  VGA_l06_g13583 : NR2D0BWP7T port map(A1 => VGA_l06_n_224, A2 => VGA_l06_n_168, ZN => VGA_l06_n_242);
  VGA_l06_g13584 : NR4D0BWP7T port map(A1 => VGA_l06_n_217, A2 => VGA_l06_n_214, A3 => VGA_l06_n_174, A4 => VGA_l06_n_104, ZN => VGA_l06_n_241);
  VGA_l06_g13585 : NR2D0BWP7T port map(A1 => VGA_l06_n_224, A2 => VGA_l06_n_139, ZN => VGA_l06_n_240);
  VGA_l06_g13586 : AOI211D0BWP7T port map(A1 => VGA_l06_n_81, A2 => VGA_l06_n_69, B => VGA_l06_n_218, C => VGA_l06_n_217, ZN => VGA_l06_n_233);
  VGA_l06_g13587 : AOI21D0BWP7T port map(A1 => VGA_l06_n_168, A2 => VGA_l06_n_177, B => VGA_l06_n_224, ZN => VGA_l06_n_232);
  VGA_l06_g13588 : IOA21D0BWP7T port map(A1 => VGA_l06_n_219, A2 => VGA_l06_n_187, B => VGA_l06_n_223, ZN => VGA_l06_n_231);
  VGA_l06_g13589 : AN3D0BWP7T port map(A1 => VGA_l06_n_227, A2 => VGA_l06_n_170, A3 => VGA_l06_n_178, Z => VGA_l06_n_230);
  VGA_l06_g13590 : IND3D0BWP7T port map(A1 => VGA_l06_n_156, B1 => VGA_l06_n_97, B2 => VGA_l06_n_219, ZN => VGA_l06_n_238);
  VGA_l06_g13592 : IND3D0BWP7T port map(A1 => VGA_l06_n_149, B1 => VGA_l06_n_97, B2 => VGA_l06_n_219, ZN => VGA_l06_n_237);
  VGA_l06_g13593 : NR4D0BWP7T port map(A1 => VGA_l06_n_214, A2 => VGA_l06_n_99, A3 => VGA_l06_n_108, A4 => VGA_l06_n_60, ZN => VGA_l06_n_236);
  VGA_l06_g13594 : IND3D0BWP7T port map(A1 => VGA_l06_n_156, B1 => VGA_l06_n_97, B2 => VGA_l06_n_221, ZN => VGA_l06_n_235);
  VGA_l06_g13595 : NR3D0BWP7T port map(A1 => VGA_l06_n_229, A2 => VGA_l06_n_107, A3 => VGA_l06_n_106, ZN => VGA_l06_n_234);
  VGA_l06_g13596 : INVD1BWP7T port map(I => VGA_l06_n_227, ZN => VGA_l06_n_228);
  VGA_l06_g13597 : ND2D0BWP7T port map(A1 => VGA_l06_n_222, A2 => VGA_l06_n_216, ZN => VGA_l06_n_229);
  VGA_l06_g13598 : NR2D0BWP7T port map(A1 => VGA_l06_n_220, A2 => VGA_l06_n_217, ZN => VGA_l06_n_227);
  VGA_l06_g13599 : CKND1BWP7T port map(I => VGA_l06_n_225, ZN => VGA_l06_n_226);
  VGA_l06_g13600 : OAI31D0BWP7T port map(A1 => VGA_l06_n_138, A2 => VGA_l06_n_178, A3 => VGA_l06_n_187, B => VGA_l06_n_221, ZN => VGA_l06_n_223);
  VGA_l06_g13601 : OAI21D0BWP7T port map(A1 => VGA_l06_n_115, A2 => VGA_l06_n_86, B => VGA_l06_n_216, ZN => VGA_l06_n_225);
  VGA_l06_g13602 : ND2D0BWP7T port map(A1 => VGA_l06_n_219, A2 => VGA_l06_n_216, ZN => VGA_l06_n_224);
  VGA_l06_g13603 : CKND1BWP7T port map(I => VGA_l06_n_221, ZN => VGA_l06_n_220);
  VGA_l06_g13604 : INR2D0BWP7T port map(A1 => VGA_l06_n_104, B1 => VGA_l06_n_213, ZN => VGA_l06_n_222);
  VGA_l06_g13605 : NR2D0BWP7T port map(A1 => VGA_l06_n_213, A2 => VGA_l06_n_103, ZN => VGA_l06_n_221);
  VGA_l06_g13606 : NR2D0BWP7T port map(A1 => VGA_l06_n_214, A2 => VGA_l06_n_102, ZN => VGA_l06_n_219);
  VGA_l06_g13608 : INVD1BWP7T port map(I => VGA_l06_n_217, ZN => VGA_l06_n_216);
  VGA_l06_g13609 : IND3D0BWP7T port map(A1 => VGA_l06_n_99, B1 => VGA_l06_n_95, B2 => VGA_l06_n_210, ZN => VGA_l06_n_215);
  VGA_l06_g13610 : ND3D0BWP7T port map(A1 => VGA_l06_n_209, A2 => VGA_l06_n_60, A3 => VGA_l06_n_47, ZN => VGA_l06_n_218);
  VGA_l06_g13611 : OAI221D0BWP7T port map(A1 => VGA_l06_n_57, A2 => VGA_l06_n_38, B1 => VGA_l06_n_8, B2 => VGA_x(8), C => VGA_l06_n_212, ZN => VGA_l06_n_217);
  VGA_l06_g13612 : OAI211D0BWP7T port map(A1 => VGA_l06_n_18, A2 => VGA_l06_n_48, B => VGA_l06_n_210, C => VGA_l06_n_75, ZN => VGA_l06_n_214);
  VGA_l06_g13613 : OAI211D0BWP7T port map(A1 => VGA_l06_n_20, A2 => VGA_l06_n_49, B => VGA_l06_n_210, C => VGA_l06_n_72, ZN => VGA_l06_n_213);
  VGA_l06_g13614 : AOI221D0BWP7T port map(A1 => VGA_l06_n_204, A2 => VGA_l06_n_153, B1 => VGA_l06_n_27, B2 => VGA_l06_n_40, C => VGA_l06_n_208, ZN => VGA_l06_n_212);
  VGA_l06_g13615 : NR4D0BWP7T port map(A1 => VGA_l06_n_205, A2 => VGA_l06_n_128, A3 => VGA_l06_n_80, A4 => VGA_l06_n_84, ZN => VGA_l06_n_211);
  VGA_l06_g13616 : OAI211D0BWP7T port map(A1 => y_pos_p(5), A2 => VGA_l06_n_197, B => VGA_l06_n_196, C => VGA_l06_n_188, ZN => VGA_l06_n_210);
  VGA_l06_g13617 : AOI211D0BWP7T port map(A1 => VGA_l06_n_197, A2 => VGA_l06_n_188, B => VGA_l06_n_99, C => VGA_l06_n_49, ZN => VGA_l06_n_209);
  VGA_l06_g13618 : OAI221D0BWP7T port map(A1 => VGA_l06_n_200, A2 => VGA_l06_n_153, B1 => VGA_l06_n_40, B2 => VGA_l06_n_27, C => VGA_l06_n_111, ZN => VGA_l06_n_208);
  VGA_l06_g13619 : IND4D0BWP7T port map(A1 => VGA_l06_n_191, B1 => VGA_l06_n_0, B2 => VGA_l06_n_129, B3 => VGA_l06_n_162, ZN => VGA_l06_n_207);
  VGA_l06_g13620 : ND3D0BWP7T port map(A1 => VGA_l06_n_198, A2 => VGA_l06_n_148, A3 => VGA_l06_n_151, ZN => VGA_l06_n_206);
  VGA_l06_g13621 : ND2D0BWP7T port map(A1 => VGA_l06_n_198, A2 => VGA_l06_n_124, ZN => VGA_l06_n_205);
  VGA_l06_g13622 : OAI211D0BWP7T port map(A1 => VGA_l06_n_16, A2 => VGA_l06_n_54, B => VGA_l06_n_189, C => VGA_l06_n_122, ZN => VGA_l06_n_204);
  VGA_l06_g13623 : AOI22D0BWP7T port map(A1 => VGA_l06_n_187, A2 => VGA_l06_n_70, B1 => VGA_l06_n_175, B2 => VGA_l06_n_178, ZN => VGA_l06_n_203);
  VGA_l06_g13624 : CKND1BWP7T port map(I => VGA_l06_n_201, ZN => VGA_l06_n_202);
  VGA_l06_g13625 : NR2D0BWP7T port map(A1 => VGA_l06_n_189, A2 => VGA_l06_n_146, ZN => VGA_l06_n_200);
  VGA_l06_g13626 : IND4D0BWP7T port map(A1 => VGA_l06_n_147, B1 => VGA_l06_n_51, B2 => VGA_l06_n_82, B3 => VGA_l06_n_157, ZN => VGA_l06_n_199);
  VGA_l06_g13627 : NR3D0BWP7T port map(A1 => VGA_l06_n_161, A2 => VGA_l06_n_171, A3 => VGA_l06_n_182, ZN => VGA_l06_n_201);
  VGA_l06_g13628 : ND3D0BWP7T port map(A1 => VGA_l06_n_172, A2 => VGA_l06_n_94, A3 => y_pos_p(5), ZN => VGA_l06_n_196);
  VGA_l06_g13629 : IND4D0BWP7T port map(A1 => VGA_l06_n_171, B1 => VGA_l06_n_82, B2 => VGA_l06_n_77, B3 => VGA_l06_n_162, ZN => VGA_l06_n_195);
  VGA_l06_g13630 : AOI21D0BWP7T port map(A1 => VGA_l06_n_31, A2 => VGA_l06_n_33, B => VGA_l06_n_194, ZN => VGA_l06_n_198);
  VGA_l06_g13631 : ND3D0BWP7T port map(A1 => VGA_l06_n_172, A2 => VGA_l06_n_52, A3 => VGA_y(5), ZN => VGA_l06_n_197);
  VGA_l06_g13632 : ND2D0BWP7T port map(A1 => VGA_l06_n_180, A2 => VGA_l06_n_142, ZN => VGA_l06_n_194);
  VGA_l06_g13633 : NR2D0BWP7T port map(A1 => VGA_l06_n_170, A2 => VGA_l06_n_171, ZN => VGA_l06_n_193);
  VGA_l06_g13634 : ND2D0BWP7T port map(A1 => VGA_l06_n_184, A2 => VGA_l06_n_71, ZN => VGA_l06_n_192);
  VGA_l06_g13635 : ND2D0BWP7T port map(A1 => VGA_l06_n_180, A2 => VGA_l06_n_116, ZN => VGA_l06_n_191);
  VGA_l06_g13636 : IND2D0BWP7T port map(A1 => VGA_l06_n_176, B1 => VGA_l06_n_51, ZN => VGA_l06_n_190);
  VGA_l06_g13637 : IND3D0BWP7T port map(A1 => VGA_l06_n_90, B1 => VGA_l06_n_51, B2 => VGA_l06_n_151, ZN => VGA_l06_n_186);
  VGA_l06_g13638 : AOI21D0BWP7T port map(A1 => VGA_l06_n_66, A2 => VGA_l06_n_30, B => VGA_l06_n_176, ZN => VGA_l06_n_185);
  VGA_l06_g13639 : AOI21D0BWP7T port map(A1 => VGA_l06_n_58, A2 => VGA_l06_n_41, B => VGA_l06_n_167, ZN => VGA_l06_n_189);
  VGA_l06_g13640 : IND3D0BWP7T port map(A1 => VGA_y(5), B1 => VGA_l06_n_94, B2 => VGA_l06_n_172, ZN => VGA_l06_n_188);
  VGA_l06_g13641 : ND2D0BWP7T port map(A1 => VGA_l06_n_169, A2 => VGA_l06_n_179, ZN => VGA_l06_n_187);
  VGA_l06_g13642 : INVD0BWP7T port map(I => VGA_l06_n_177, ZN => VGA_l06_n_178);
  VGA_l06_g13643 : IND2D0BWP7T port map(A1 => VGA_l06_n_86, B1 => VGA_l06_n_148, ZN => VGA_l06_n_175);
  VGA_l06_g13644 : INR2D0BWP7T port map(A1 => VGA_l06_n_148, B1 => VGA_l06_n_70, ZN => VGA_l06_n_184);
  VGA_l06_g13645 : IND2D0BWP7T port map(A1 => VGA_l06_n_147, B1 => VGA_l06_n_71, ZN => VGA_l06_n_183);
  VGA_l06_g13646 : IND2D0BWP7T port map(A1 => VGA_l06_n_91, B1 => VGA_l06_n_164, ZN => VGA_l06_n_182);
  VGA_l06_g13647 : IND2D0BWP7T port map(A1 => VGA_l06_n_117, B1 => VGA_l06_n_148, ZN => VGA_l06_n_181);
  VGA_l06_g13648 : INR2D0BWP7T port map(A1 => VGA_l06_n_157, B1 => VGA_l06_n_117, ZN => VGA_l06_n_180);
  VGA_l06_g13649 : IND2D0BWP7T port map(A1 => VGA_l06_n_163, B1 => VGA_l06_n_96, ZN => VGA_l06_n_179);
  VGA_l06_g13650 : ND2D0BWP7T port map(A1 => VGA_l06_n_4, A2 => VGA_l06_n_97, ZN => VGA_l06_n_177);
  VGA_l06_g13651 : ND2D0BWP7T port map(A1 => VGA_l06_n_157, A2 => VGA_l06_n_136, ZN => VGA_l06_n_176);
  VGA_l06_g13652 : OA221D0BWP7T port map(A1 => VGA_l06_n_113, A2 => VGA_l06_n_73, B1 => VGA_l06_n_41, B2 => VGA_l06_n_58, C => VGA_l06_n_74, Z => VGA_l06_n_167);
  VGA_l06_g13653 : IND4D0BWP7T port map(A1 => VGA_l06_n_92, B1 => VGA_l06_n_78, B2 => VGA_l06_n_123, B3 => VGA_l06_n_142, ZN => VGA_l06_n_166);
  VGA_l06_g13654 : OAI21D0BWP7T port map(A1 => VGA_l06_n_63, A2 => VGA_l06_n_29, B => VGA_l06_n_150, ZN => VGA_l06_n_165);
  VGA_l06_g13655 : IND2D0BWP7T port map(A1 => VGA_l06_n_96, B1 => VGA_l06_n_152, ZN => VGA_l06_n_174);
  VGA_l06_g13656 : AO211D0BWP7T port map(A1 => VGA_l06_n_67, A2 => VGA_l06_n_15, B => VGA_l06_n_147, C => VGA_l06_n_132, Z => VGA_l06_n_173);
  VGA_l06_g13657 : AOI211D0BWP7T port map(A1 => VGA_l06_n_55, A2 => VGA_l06_n_24, B => VGA_l06_n_145, C => VGA_l06_n_114, ZN => VGA_l06_n_172);
  VGA_l06_g13658 : OAI21D0BWP7T port map(A1 => VGA_l06_n_89, A2 => VGA_l06_n_29, B => VGA_l06_n_150, ZN => VGA_l06_n_171);
  VGA_l06_g13659 : OAI21D0BWP7T port map(A1 => VGA_l06_n_118, A2 => VGA_l06_n_12, B => VGA_l06_n_160, ZN => VGA_l06_n_170);
  VGA_l06_g13660 : IND2D0BWP7T port map(A1 => VGA_l06_n_1, B1 => VGA_l06_n_96, ZN => VGA_l06_n_169);
  VGA_l06_g13661 : ND2D0BWP7T port map(A1 => VGA_l06_n_152, A2 => VGA_l06_n_96, ZN => VGA_l06_n_168);
  VGA_l06_g13662 : CKND1BWP7T port map(I => VGA_l06_n_160, ZN => VGA_l06_n_161);
  VGA_l06_g13663 : CKND1BWP7T port map(I => VGA_l06_n_158, ZN => VGA_l06_n_159);
  VGA_l06_g13664 : CKND1BWP7T port map(I => VGA_l06_n_3, ZN => VGA_l06_n_155);
  VGA_l06_g13665 : INR2D0BWP7T port map(A1 => VGA_l06_n_140, B1 => VGA_l06_n_84, ZN => VGA_l06_n_164);
  VGA_l06_g13666 : ND2D0BWP7T port map(A1 => VGA_l06_n_2, A2 => VGA_l06_n_105, ZN => VGA_l06_n_163);
  VGA_l06_g13668 : NR2D0BWP7T port map(A1 => VGA_l06_n_133, A2 => VGA_l06_n_132, ZN => VGA_l06_n_162);
  VGA_l06_g13669 : NR2D0BWP7T port map(A1 => VGA_l06_n_137, A2 => VGA_l06_n_76, ZN => VGA_l06_n_160);
  VGA_l06_g13670 : ND2D0BWP7T port map(A1 => VGA_l06_n_129, A2 => VGA_l06_n_32, ZN => VGA_l06_n_158);
  VGA_l06_g13671 : NR2D0BWP7T port map(A1 => VGA_l06_n_143, A2 => VGA_l06_n_92, ZN => VGA_l06_n_157);
  VGA_l06_g13672 : ND2D0BWP7T port map(A1 => VGA_l06_n_141, A2 => VGA_l06_n_109, ZN => VGA_l06_n_156);
  VGA_l06_g13674 : ND2D0BWP7T port map(A1 => VGA_l06_n_136, A2 => VGA_l06_n_119, ZN => VGA_l06_n_154);
  VGA_l06_g13675 : OAI31D0BWP7T port map(A1 => VGA_l06_n_7, A2 => VGA_x(5), A3 => VGA_l06_n_53, B => VGA_l06_n_112, ZN => VGA_l06_n_146);
  VGA_l06_g13676 : OAI221D0BWP7T port map(A1 => VGA_l06_n_56, A2 => VGA_l06_n_43, B1 => VGA_y(9), B2 => VGA_l06_n_42, C => VGA_l06_n_125, ZN => VGA_l06_n_145);
  VGA_l06_g13677 : OAI21D0BWP7T port map(A1 => VGA_l06_n_118, A2 => VGA_l06_n_32, B => VGA_l06_n_131, ZN => VGA_l06_n_144);
  VGA_l06_g13678 : ND2D0BWP7T port map(A1 => VGA_l06_n_127, A2 => VGA_l06_n_122, ZN => VGA_l06_n_153);
  VGA_l06_g13680 : INR2D0BWP7T port map(A1 => VGA_l06_n_141, B1 => VGA_l06_n_109, ZN => VGA_l06_n_152);
  VGA_l06_g13681 : IAO21D0BWP7T port map(A1 => VGA_l06_n_89, A2 => VGA_l06_n_32, B => VGA_l06_n_128, ZN => VGA_l06_n_151);
  VGA_l06_g13682 : AOI211D0BWP7T port map(A1 => VGA_l06_n_85, A2 => VGA_l06_n_30, B => VGA_l06_n_87, C => VGA_l06_n_79, ZN => VGA_l06_n_150);
  VGA_l06_g13683 : ND3D0BWP7T port map(A1 => VGA_l06_n_100, A2 => VGA_l06_n_62, A3 => VGA_l06_n_50, ZN => VGA_l06_n_149);
  VGA_l06_g13684 : AOI211D0BWP7T port map(A1 => VGA_l06_n_61, A2 => VGA_l06_n_13, B => VGA_l06_n_115, C => VGA_l06_n_84, ZN => VGA_l06_n_148);
  VGA_l06_g13685 : AO21D0BWP7T port map(A1 => VGA_l06_n_61, A2 => VGA_l06_n_15, B => VGA_l06_n_133, Z => VGA_l06_n_147);
  VGA_l06_g13687 : CKND1BWP7T port map(I => VGA_l06_n_139, ZN => VGA_l06_n_138);
  VGA_l06_g13688 : INVD0BWP7T port map(I => VGA_l06_n_136, ZN => VGA_l06_n_135);
  VGA_l06_g13689 : IND2D0BWP7T port map(A1 => VGA_l06_n_99, B1 => VGA_l06_n_108, ZN => VGA_l06_n_134);
  VGA_l06_g13690 : IND2D0BWP7T port map(A1 => VGA_l06_n_79, B1 => VGA_l06_n_119, ZN => VGA_l06_n_143);
  VGA_l06_g13691 : INR2D0BWP7T port map(A1 => VGA_l06_n_51, B1 => VGA_l06_n_121, ZN => VGA_l06_n_142);
  VGA_l06_g13692 : NR2D0BWP7T port map(A1 => VGA_l06_n_101, A2 => VGA_l06_n_50, ZN => VGA_l06_n_141);
  VGA_l06_g13693 : OA21D0BWP7T port map(A1 => VGA_l06_n_88, A2 => VGA_l06_n_12, B => VGA_l06_n_81, Z => VGA_l06_n_140);
  VGA_l06_g13695 : IND2D0BWP7T port map(A1 => VGA_l06_n_106, B1 => VGA_l06_n_107, ZN => VGA_l06_n_139);
  VGA_l06_g13696 : OR2D0BWP7T port map(A1 => VGA_l06_n_117, A2 => VGA_l06_n_80, Z => VGA_l06_n_137);
  VGA_l06_g13697 : NR2D0BWP7T port map(A1 => VGA_l06_n_115, A2 => VGA_l06_n_117, ZN => VGA_l06_n_136);
  VGA_l06_g13698 : CKND1BWP7T port map(I => VGA_l06_n_130, ZN => VGA_l06_n_131);
  VGA_l06_g13699 : MOAI22D0BWP7T port map(A1 => VGA_l06_n_53, A2 => VGA_l06_n_26, B1 => VGA_l06_n_54, B2 => VGA_l06_n_16, ZN => VGA_l06_n_127);
  VGA_l06_g13700 : AOI21D0BWP7T port map(A1 => VGA_l06_n_93, A2 => VGA_l06_n_13, B => VGA_l06_n_84, ZN => VGA_l06_n_126);
  VGA_l06_g13701 : AOI22D0BWP7T port map(A1 => VGA_l06_n_56, A2 => VGA_l06_n_43, B1 => VGA_l06_n_42, B2 => VGA_y(9), ZN => VGA_l06_n_125);
  VGA_l06_g13702 : IOA21D0BWP7T port map(A1 => VGA_l06_n_89, A2 => VGA_l06_n_64, B => VGA_l06_n_31, ZN => VGA_l06_n_124);
  VGA_l06_g13703 : OAI21D0BWP7T port map(A1 => VGA_l06_n_63, A2 => VGA_l06_n_14, B => VGA_l06_n_120, ZN => VGA_l06_n_133);
  VGA_l06_g13704 : IND3D0BWP7T port map(A1 => VGA_l06_n_84, B1 => VGA_l06_n_81, B2 => VGA_l06_n_78, ZN => VGA_l06_n_132);
  VGA_l06_g13705 : IND3D0BWP7T port map(A1 => VGA_l06_n_84, B1 => VGA_l06_n_51, B2 => VGA_l06_n_78, ZN => VGA_l06_n_130);
  VGA_l06_g13706 : IAO21D0BWP7T port map(A1 => VGA_l06_n_88, A2 => VGA_l06_n_32, B => VGA_l06_n_83, ZN => VGA_l06_n_129);
  VGA_l06_g13707 : IAO21D0BWP7T port map(A1 => VGA_l06_n_85, A2 => VGA_l06_n_61, B => VGA_l06_n_32, ZN => VGA_l06_n_128);
  VGA_l06_g13709 : INVD0BWP7T port map(I => VGA_l06_n_116, ZN => VGA_l06_n_115);
  VGA_l06_g13710 : NR2D0BWP7T port map(A1 => VGA_l06_n_55, A2 => VGA_l06_n_24, ZN => VGA_l06_n_114);
  VGA_l06_g13711 : MOAI22D0BWP7T port map(A1 => VGA_l06_n_11, A2 => x_pos_p(1), B1 => VGA_l06_n_44, B2 => VGA_x(0), ZN => VGA_l06_n_113);
  VGA_l06_g13712 : IND2D0BWP7T port map(A1 => VGA_l06_n_54, B1 => VGA_l06_n_16, ZN => VGA_l06_n_112);
  VGA_l06_g13713 : ND2D0BWP7T port map(A1 => VGA_l06_n_57, A2 => VGA_l06_n_38, ZN => VGA_l06_n_111);
  VGA_l06_g13714 : AOI21D0BWP7T port map(A1 => VGA_l06_n_63, A2 => VGA_l06_n_65, B => VGA_l06_n_32, ZN => VGA_l06_n_110);
  VGA_l06_g13715 : ND2D0BWP7T port map(A1 => VGA_l06_n_85, A2 => VGA_l06_n_13, ZN => VGA_l06_n_123);
  VGA_l06_g13716 : ND2D0BWP7T port map(A1 => VGA_l06_n_53, A2 => VGA_l06_n_26, ZN => VGA_l06_n_122);
  VGA_l06_g13717 : OR2D0BWP7T port map(A1 => VGA_l06_n_90, A2 => VGA_l06_n_83, Z => VGA_l06_n_121);
  VGA_l06_g13718 : ND2D0BWP7T port map(A1 => VGA_l06_n_85, A2 => VGA_l06_n_15, ZN => VGA_l06_n_120);
  VGA_l06_g13719 : NR2D0BWP7T port map(A1 => VGA_l06_n_76, A2 => VGA_l06_n_87, ZN => VGA_l06_n_119);
  VGA_l06_g13720 : NR2D0BWP7T port map(A1 => VGA_l06_n_85, A2 => VGA_l06_n_93, ZN => VGA_l06_n_118);
  VGA_l06_g13721 : IND2D0BWP7T port map(A1 => VGA_l06_n_86, B1 => VGA_l06_n_82, ZN => VGA_l06_n_117);
  VGA_l06_g13722 : NR2D0BWP7T port map(A1 => VGA_l06_n_80, A2 => VGA_l06_n_91, ZN => VGA_l06_n_116);
  VGA_l06_g13723 : CKND1BWP7T port map(I => VGA_l06_n_102, ZN => VGA_l06_n_103);
  VGA_l06_g13726 : CKND1BWP7T port map(I => VGA_l06_n_97, ZN => VGA_l06_n_98);
  VGA_l06_g13727 : MAOI22D0BWP7T port map(A1 => VGA_l06_n_49, A2 => VGA_y(4), B1 => VGA_l06_n_49, B2 => VGA_y(4), ZN => VGA_l06_n_95);
  VGA_l06_g13728 : MOAI22D0BWP7T port map(A1 => VGA_l06_n_46, A2 => VGA_l06_n_34, B1 => VGA_l06_n_46, B2 => VGA_l06_n_34, ZN => VGA_l06_n_109);
  VGA_l06_g13729 : MOAI22D0BWP7T port map(A1 => VGA_l06_n_47, A2 => VGA_y(3), B1 => VGA_l06_n_47, B2 => VGA_y(3), ZN => VGA_l06_n_108);
  VGA_l06_g13730 : MAOI22D0BWP7T port map(A1 => VGA_l06_n_59, A2 => VGA_y(2), B1 => VGA_l06_n_59, B2 => VGA_y(2), ZN => VGA_l06_n_107);
  VGA_l06_g13731 : IND3D0BWP7T port map(A1 => VGA_l06_n_62, B1 => VGA_l06_n_50, B2 => VGA_l06_n_46, ZN => VGA_l06_n_106);
  VGA_l06_g13732 : MOAI22D0BWP7T port map(A1 => VGA_l06_n_46, A2 => VGA_l06_n_19, B1 => VGA_l06_n_46, B2 => VGA_l06_n_19, ZN => VGA_l06_n_105);
  VGA_l06_g13733 : MOAI22D0BWP7T port map(A1 => VGA_l06_n_47, A2 => VGA_l06_n_37, B1 => VGA_l06_n_47, B2 => VGA_l06_n_37, ZN => VGA_l06_n_104);
  VGA_l06_g13734 : MOAI22D0BWP7T port map(A1 => VGA_l06_n_47, A2 => VGA_l06_n_35, B1 => VGA_l06_n_47, B2 => VGA_l06_n_35, ZN => VGA_l06_n_102);
  VGA_l06_g13735 : MOAI22D0BWP7T port map(A1 => VGA_l06_n_62, A2 => VGA_y(0), B1 => VGA_l06_n_62, B2 => VGA_y(0), ZN => VGA_l06_n_101);
  VGA_l06_g13736 : MOAI22D0BWP7T port map(A1 => VGA_l06_n_46, A2 => VGA_y(1), B1 => VGA_l06_n_46, B2 => VGA_y(1), ZN => VGA_l06_n_100);
  VGA_l06_g13737 : IND3D0BWP7T port map(A1 => VGA_l06_n_62, B1 => VGA_l06_n_50, B2 => VGA_l06_n_45, ZN => VGA_l06_n_99);
  VGA_l06_g13738 : MOAI22D0BWP7T port map(A1 => VGA_l06_n_59, A2 => VGA_l06_n_36, B1 => VGA_l06_n_59, B2 => VGA_l06_n_36, ZN => VGA_l06_n_97);
  VGA_l06_g13739 : MOAI22D0BWP7T port map(A1 => VGA_l06_n_59, A2 => VGA_l06_n_23, B1 => VGA_l06_n_59, B2 => VGA_l06_n_23, ZN => VGA_l06_n_96);
  VGA_l06_g13740 : CKND1BWP7T port map(I => VGA_l06_n_52, ZN => VGA_l06_n_94);
  VGA_l06_g13741 : OR2D0BWP7T port map(A1 => VGA_l06_n_67, A2 => VGA_l06_n_61, Z => VGA_l06_n_93);
  VGA_l06_g13742 : NR2D0BWP7T port map(A1 => VGA_l06_n_0, A2 => VGA_l06_n_29, ZN => VGA_l06_n_92);
  VGA_l06_g13743 : INR2D0BWP7T port map(A1 => VGA_l06_n_66, B1 => VGA_l06_n_12, ZN => VGA_l06_n_91);
  VGA_l06_g13744 : INR2D0BWP7T port map(A1 => VGA_l06_n_68, B1 => VGA_l06_n_29, ZN => VGA_l06_n_90);
  VGA_l06_g13745 : INR2D0BWP7T port map(A1 => VGA_l06_n_63, B1 => VGA_l06_n_68, ZN => VGA_l06_n_89);
  VGA_l06_g13746 : NR2D0BWP7T port map(A1 => VGA_l06_n_61, A2 => VGA_l06_n_33, ZN => VGA_l06_n_88);
  VGA_l06_g13747 : INR2D0BWP7T port map(A1 => VGA_l06_n_67, B1 => VGA_l06_n_29, ZN => VGA_l06_n_87);
  VGA_l06_g13748 : INR2D0BWP7T port map(A1 => VGA_l06_n_68, B1 => VGA_l06_n_12, ZN => VGA_l06_n_86);
  VGA_l06_g13749 : IND2D0BWP7T port map(A1 => VGA_l06_n_66, B1 => VGA_l06_n_0, ZN => VGA_l06_n_85);
  VGA_l06_g13750 : NR2D0BWP7T port map(A1 => VGA_l06_n_0, A2 => VGA_l06_n_12, ZN => VGA_l06_n_84);
  VGA_l06_g13751 : CKND1BWP7T port map(I => VGA_l06_n_76, ZN => VGA_l06_n_77);
  VGA_l06_g13752 : ND2D0BWP7T port map(A1 => VGA_l06_n_48, A2 => VGA_l06_n_18, ZN => VGA_l06_n_75);
  VGA_l06_g13753 : OAI22D0BWP7T port map(A1 => VGA_l06_n_39, A2 => VGA_l06_n_25, B1 => VGA_l06_n_10, B2 => x_pos_p(2), ZN => VGA_l06_n_74);
  VGA_l06_g13754 : AOI211D0BWP7T port map(A1 => VGA_l06_n_10, A2 => x_pos_p(2), B => VGA_l06_n_39, C => VGA_l06_n_25, ZN => VGA_l06_n_73);
  VGA_l06_g13755 : ND2D0BWP7T port map(A1 => VGA_l06_n_49, A2 => VGA_l06_n_20, ZN => VGA_l06_n_72);
  VGA_l06_g13756 : NR2D0BWP7T port map(A1 => VGA_l06_n_64, A2 => VGA_l06_n_29, ZN => VGA_l06_n_83);
  VGA_l06_g13757 : IND2D0BWP7T port map(A1 => VGA_l06_n_64, B1 => VGA_l06_n_13, ZN => VGA_l06_n_82);
  VGA_l06_g13758 : IND2D0BWP7T port map(A1 => VGA_l06_n_64, B1 => VGA_l06_n_15, ZN => VGA_l06_n_81);
  VGA_l06_g13759 : NR2D0BWP7T port map(A1 => VGA_l06_n_63, A2 => VGA_l06_n_12, ZN => VGA_l06_n_80);
  VGA_l06_g13760 : INR2D0BWP7T port map(A1 => VGA_l06_n_61, B1 => VGA_l06_n_29, ZN => VGA_l06_n_79);
  VGA_l06_g13761 : IND2D0BWP7T port map(A1 => VGA_l06_n_65, B1 => VGA_l06_n_13, ZN => VGA_l06_n_78);
  VGA_l06_g13762 : NR2D0BWP7T port map(A1 => VGA_l06_n_65, A2 => VGA_l06_n_29, ZN => VGA_l06_n_76);
  VGA_l06_g13763 : CKND1BWP7T port map(I => VGA_l06_n_69, ZN => VGA_l06_n_70);
  VGA_l06_g13764 : INVD1BWP7T port map(I => VGA_l06_n_60, ZN => VGA_l06_n_59);
  VGA_l06_g13765 : IND2D0BWP7T port map(A1 => VGA_l06_n_17, B1 => VGA_l06_n_15, ZN => VGA_l06_n_71);
  VGA_l06_g13766 : ND2D0BWP7T port map(A1 => VGA_l06_n_13, A2 => VGA_l06_n_33, ZN => VGA_l06_n_69);
  VGA_l06_g13767 : NR2D0BWP7T port map(A1 => VGA_l06_n_17, A2 => VGA_draw_count4(0), ZN => VGA_l06_n_68);
  VGA_l06_g13768 : AN2D1BWP7T port map(A1 => VGA_l06_n_33, A2 => VGA_draw_count4(0), Z => VGA_l06_n_67);
  VGA_l06_g13769 : NR2D0BWP7T port map(A1 => VGA_l06_n_21, A2 => VGA_draw_count4(0), ZN => VGA_l06_n_66);
  VGA_l06_g13770 : IND2D0BWP7T port map(A1 => VGA_draw_count4(0), B1 => VGA_l06_n_33, ZN => VGA_l06_n_65);
  VGA_l06_g13772 : IND2D0BWP7T port map(A1 => VGA_l06_n_17, B1 => VGA_draw_count4(0), ZN => VGA_l06_n_64);
  VGA_l06_g13773 : ND2D0BWP7T port map(A1 => VGA_l06_n_22, A2 => VGA_draw_count4(0), ZN => VGA_l06_n_63);
  VGA_l06_g13774 : ND2D0BWP7T port map(A1 => VGA_l06_n_34, A2 => VGA_l06_n_19, ZN => VGA_l06_n_62);
  VGA_l06_g13775 : NR2D0BWP7T port map(A1 => VGA_l06_n_28, A2 => VGA_draw_count4(0), ZN => VGA_l06_n_61);
  VGA_l06_g13776 : INR2D0BWP7T port map(A1 => VGA_l06_n_35, B1 => VGA_l06_n_37, ZN => VGA_l06_n_60);
  VGA_l06_g13777 : CKND1BWP7T port map(I => VGA_l06_n_49, ZN => VGA_l06_n_48);
  VGA_l06_g13778 : INVD1BWP7T port map(I => VGA_l06_n_45, ZN => VGA_l06_n_46);
  VGA_l06_g13779 : AOI21D0BWP7T port map(A1 => VGA_l06_n_11, A2 => x_pos_p(1), B => x_pos_p(0), ZN => VGA_l06_n_44);
  VGA_l06_g13780 : AO21D0BWP7T port map(A1 => VGA_x(4), A2 => VGA_l06_n_9, B => VGA_l06_n_16, Z => VGA_l06_n_58);
  VGA_l06_g13781 : MAOI22D0BWP7T port map(A1 => VGA_x(7), A2 => x_pos_p(7), B1 => VGA_x(7), B2 => x_pos_p(7), ZN => VGA_l06_n_57);
  VGA_l06_g13782 : MAOI22D0BWP7T port map(A1 => VGA_y(7), A2 => y_pos_p(7), B1 => VGA_y(7), B2 => y_pos_p(7), ZN => VGA_l06_n_56);
  VGA_l06_g13783 : MAOI22D0BWP7T port map(A1 => VGA_y(8), A2 => y_pos_p(8), B1 => VGA_y(8), B2 => y_pos_p(8), ZN => VGA_l06_n_55);
  VGA_l06_g13784 : MAOI22D0BWP7T port map(A1 => VGA_x(5), A2 => x_pos_p(5), B1 => VGA_x(5), B2 => x_pos_p(5), ZN => VGA_l06_n_54);
  VGA_l06_g13785 : MOAI22D0BWP7T port map(A1 => VGA_x(6), A2 => x_pos_p(6), B1 => VGA_x(6), B2 => x_pos_p(6), ZN => VGA_l06_n_53);
  VGA_l06_g13786 : MOAI22D0BWP7T port map(A1 => VGA_y(6), A2 => y_pos_p(6), B1 => VGA_y(6), B2 => y_pos_p(6), ZN => VGA_l06_n_52);
  VGA_l06_g13787 : ND2D0BWP7T port map(A1 => VGA_l06_n_30, A2 => VGA_l06_n_22, ZN => VGA_l06_n_51);
  VGA_l06_g13788 : XNR2D1BWP7T port map(A1 => VGA_y(0), A2 => y_pos_p(0), ZN => VGA_l06_n_50);
  VGA_l06_g13789 : MOAI22D0BWP7T port map(A1 => VGA_y(5), A2 => y_pos_p(5), B1 => VGA_y(5), B2 => y_pos_p(5), ZN => VGA_l06_n_49);
  VGA_l06_g13790 : AN2D1BWP7T port map(A1 => VGA_l06_n_20, A2 => VGA_l06_n_18, Z => VGA_l06_n_47);
  VGA_l06_g13791 : INR2D0BWP7T port map(A1 => VGA_l06_n_36, B1 => VGA_l06_n_23, ZN => VGA_l06_n_45);
  VGA_l06_g13792 : INVD0BWP7T port map(I => VGA_l06_n_32, ZN => VGA_l06_n_31);
  VGA_l06_g13793 : INVD1BWP7T port map(I => VGA_l06_n_30, ZN => VGA_l06_n_29);
  VGA_l06_g13794 : IND2D0BWP7T port map(A1 => VGA_y(6), B1 => y_pos_p(6), ZN => VGA_l06_n_43);
  VGA_l06_g13795 : IND2D0BWP7T port map(A1 => VGA_y(8), B1 => y_pos_p(8), ZN => VGA_l06_n_42);
  VGA_l06_g13796 : IND2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_p(3), ZN => VGA_l06_n_41);
  VGA_l06_g13797 : INR2D0BWP7T port map(A1 => VGA_x(8), B1 => x_pos_p(8), ZN => VGA_l06_n_40);
  VGA_l06_g13798 : AN2D1BWP7T port map(A1 => VGA_x(3), A2 => x_pos_p(3), Z => VGA_l06_n_39);
  VGA_l06_g13799 : INR2D0BWP7T port map(A1 => VGA_x(6), B1 => x_pos_p(6), ZN => VGA_l06_n_38);
  VGA_l06_g13800 : INR2D0BWP7T port map(A1 => VGA_y(3), B1 => y_pos_p(3), ZN => VGA_l06_n_37);
  VGA_l06_g13801 : IND2D0BWP7T port map(A1 => y_pos_p(2), B1 => VGA_y(2), ZN => VGA_l06_n_36);
  VGA_l06_g13802 : IND2D0BWP7T port map(A1 => VGA_y(3), B1 => y_pos_p(3), ZN => VGA_l06_n_35);
  VGA_l06_g13803 : IND2D0BWP7T port map(A1 => VGA_y(1), B1 => y_pos_p(1), ZN => VGA_l06_n_34);
  VGA_l06_g13804 : NR2D0BWP7T port map(A1 => VGA_draw_count4(2), A2 => VGA_draw_count4(1), ZN => VGA_l06_n_33);
  VGA_l06_g13805 : ND2D0BWP7T port map(A1 => VGA_draw_count4(3), A2 => VGA_draw_count4(4), ZN => VGA_l06_n_32);
  VGA_l06_g13806 : INR2D0BWP7T port map(A1 => VGA_draw_count4(4), B1 => VGA_draw_count4(3), ZN => VGA_l06_n_30);
  VGA_l06_g13808 : CKND1BWP7T port map(I => VGA_l06_n_21, ZN => VGA_l06_n_22);
  VGA_l06_g13809 : CKND1BWP7T port map(I => VGA_l06_n_15, ZN => VGA_l06_n_14);
  VGA_l06_g13810 : INVD1BWP7T port map(I => VGA_l06_n_13, ZN => VGA_l06_n_12);
  VGA_l06_g13811 : IND2D0BWP7T port map(A1 => VGA_draw_count4(2), B1 => VGA_draw_count4(1), ZN => VGA_l06_n_28);
  VGA_l06_g13812 : IND2D0BWP7T port map(A1 => VGA_x(7), B1 => x_pos_p(7), ZN => VGA_l06_n_27);
  VGA_l06_g13813 : INR2D0BWP7T port map(A1 => VGA_x(5), B1 => x_pos_p(5), ZN => VGA_l06_n_26);
  VGA_l06_g13814 : NR2D0BWP7T port map(A1 => VGA_x(3), A2 => x_pos_p(3), ZN => VGA_l06_n_25);
  VGA_l06_g13815 : IND2D0BWP7T port map(A1 => VGA_y(7), B1 => y_pos_p(7), ZN => VGA_l06_n_24);
  VGA_l06_g13816 : INR2D0BWP7T port map(A1 => y_pos_p(2), B1 => VGA_y(2), ZN => VGA_l06_n_23);
  VGA_l06_g13817 : IND2D0BWP7T port map(A1 => VGA_draw_count4(1), B1 => VGA_draw_count4(2), ZN => VGA_l06_n_21);
  VGA_l06_g13818 : IND2D0BWP7T port map(A1 => VGA_y(4), B1 => y_pos_p(4), ZN => VGA_l06_n_20);
  VGA_l06_g13819 : IND2D0BWP7T port map(A1 => y_pos_p(1), B1 => VGA_y(1), ZN => VGA_l06_n_19);
  VGA_l06_g13820 : IND2D0BWP7T port map(A1 => y_pos_p(4), B1 => VGA_y(4), ZN => VGA_l06_n_18);
  VGA_l06_g13821 : ND2D0BWP7T port map(A1 => VGA_draw_count4(1), A2 => VGA_draw_count4(2), ZN => VGA_l06_n_17);
  VGA_l06_g13822 : NR2D0BWP7T port map(A1 => VGA_x(4), A2 => VGA_l06_n_9, ZN => VGA_l06_n_16);
  VGA_l06_g13823 : NR2D0BWP7T port map(A1 => VGA_draw_count4(4), A2 => VGA_draw_count4(3), ZN => VGA_l06_n_15);
  VGA_l06_g13824 : INR2D0BWP7T port map(A1 => VGA_draw_count4(3), B1 => VGA_draw_count4(4), ZN => VGA_l06_n_13);
  VGA_l06_g13825 : CKND1BWP7T port map(I => VGA_x(1), ZN => VGA_l06_n_11);
  VGA_l06_g13826 : CKND1BWP7T port map(I => VGA_x(2), ZN => VGA_l06_n_10);
  VGA_l06_g13827 : CKND1BWP7T port map(I => x_pos_p(4), ZN => VGA_l06_n_9);
  VGA_l06_g13828 : CKND1BWP7T port map(I => x_pos_p(8), ZN => VGA_l06_n_8);
  VGA_l06_g13829 : CKND1BWP7T port map(I => x_pos_p(5), ZN => VGA_l06_n_7);
  VGA_l06_g2 : IND2D1BWP7T port map(A1 => VGA_l06_n_247, B1 => VGA_l06_n_4, ZN => VGA_l06_n_6);
  VGA_l06_g13830 : OA21D0BWP7T port map(A1 => VGA_l06_n_220, A2 => VGA_l06_n_168, B => VGA_l06_n_218, Z => VGA_l06_n_5);
  VGA_l06_g13831 : INR2D1BWP7T port map(A1 => VGA_l06_n_2, B1 => VGA_l06_n_105, ZN => VGA_l06_n_4);
  VGA_l06_g13832 : INR2D1BWP7T port map(A1 => VGA_l06_n_119, B1 => VGA_l06_n_137, ZN => VGA_l06_n_3);
  VGA_l06_g13833 : INR2D1BWP7T port map(A1 => VGA_l06_n_101, B1 => VGA_l06_n_50, ZN => VGA_l06_n_2);
  VGA_l06_g13834 : IND3D1BWP7T port map(A1 => VGA_l06_n_100, B1 => VGA_l06_n_62, B2 => VGA_l06_n_50, ZN => VGA_l06_n_1);
  VGA_l06_g13835 : IND2D1BWP7T port map(A1 => VGA_l06_n_28, B1 => VGA_draw_count4(0), ZN => VGA_l06_n_0);
  VGA_l042_count_reg_2 : DFCNQD1BWP7T port map(CDN => VGA_l042_n_0, CP => clk, D => VGA_l042_n_6, Q => VGA_draw_count2(2));
  VGA_l042_g59 : INR2D0BWP7T port map(A1 => VGA_enable2, B1 => VGA_l042_n_5, ZN => VGA_l042_n_6);
  VGA_l042_count_reg_1 : DFCNQD1BWP7T port map(CDN => VGA_l042_n_0, CP => clk, D => VGA_l042_n_4, Q => VGA_draw_count2(1));
  VGA_l042_g61 : MAOI22D0BWP7T port map(A1 => VGA_l042_n_1, A2 => VGA_draw_count2(2), B1 => VGA_l042_n_1, B2 => VGA_draw_count2(2), ZN => VGA_l042_n_5);
  VGA_l042_g62 : INR2D0BWP7T port map(A1 => VGA_enable2, B1 => VGA_l042_n_3, ZN => VGA_l042_n_4);
  VGA_l042_count_reg_0 : DFCNQD1BWP7T port map(CDN => VGA_l042_n_0, CP => clk, D => VGA_l042_n_2, Q => VGA_draw_count2(0));
  VGA_l042_g64 : XNR2D1BWP7T port map(A1 => VGA_draw_count2(0), A2 => VGA_draw_count2(1), ZN => VGA_l042_n_3);
  VGA_l042_g65 : INR2D0BWP7T port map(A1 => VGA_enable2, B1 => VGA_draw_count2(0), ZN => VGA_l042_n_2);
  VGA_l042_g66 : ND2D0BWP7T port map(A1 => VGA_draw_count2(0), A2 => VGA_draw_count2(1), ZN => VGA_l042_n_1);
  VGA_l042_g67 : INVD0BWP7T port map(I => reset, ZN => VGA_l042_n_0);
  VGA_l043_count_reg_2 : DFCNQD1BWP7T port map(CDN => VGA_l043_n_0, CP => clk, D => VGA_l043_n_6, Q => VGA_draw_count3(2));
  VGA_l043_g59 : INR2D0BWP7T port map(A1 => VGA_enable3, B1 => VGA_l043_n_5, ZN => VGA_l043_n_6);
  VGA_l043_count_reg_1 : DFCNQD1BWP7T port map(CDN => VGA_l043_n_0, CP => clk, D => VGA_l043_n_4, Q => VGA_draw_count3(1));
  VGA_l043_g61 : MAOI22D0BWP7T port map(A1 => VGA_l043_n_1, A2 => VGA_draw_count3(2), B1 => VGA_l043_n_1, B2 => VGA_draw_count3(2), ZN => VGA_l043_n_5);
  VGA_l043_g62 : INR2D0BWP7T port map(A1 => VGA_enable3, B1 => VGA_l043_n_3, ZN => VGA_l043_n_4);
  VGA_l043_count_reg_0 : DFCNQD1BWP7T port map(CDN => VGA_l043_n_0, CP => clk, D => VGA_l043_n_2, Q => VGA_draw_count3(0));
  VGA_l043_g64 : XNR2D1BWP7T port map(A1 => VGA_draw_count3(0), A2 => VGA_draw_count3(1), ZN => VGA_l043_n_3);
  VGA_l043_g65 : INR2D0BWP7T port map(A1 => VGA_enable3, B1 => VGA_draw_count3(0), ZN => VGA_l043_n_2);
  VGA_l043_g66 : ND2D0BWP7T port map(A1 => VGA_draw_count3(0), A2 => VGA_draw_count3(1), ZN => VGA_l043_n_1);
  VGA_l043_g67 : INVD0BWP7T port map(I => reset, ZN => VGA_l043_n_0);
  Enemy_spawning_rngg_g34 : XNR4D0BWP7T port map(A1 => y_e_spawn_1(0), A2 => y_e_spawn_3(1), A3 => y_e_spawn_3(3), A4 => y_e_spawn_1(7), ZN => Enemy_spawning_rngg_xor_input);
  Enemy_spawning_rngg_d10_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d10_n_0, CP => n_5, D => y_e_spawn_2(3), Q => y_e_spawn_1(3));
  Enemy_spawning_rngg_d10_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d10_n_0);
  Enemy_spawning_rngg_d11_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d11_n_0, CP => n_5, D => y_e_spawn_1(3), Q => y_e_spawn_2(1));
  Enemy_spawning_rngg_d11_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d11_n_0);
  Enemy_spawning_rngg_d12_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d12_n_0, CP => n_5, D => y_e_spawn_2(1), Q => y_e_spawn_1(2));
  Enemy_spawning_rngg_d12_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d12_n_0);
  Enemy_spawning_rngg_d13_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d13_n_0, CP => n_5, D => y_e_spawn_1(2), Q => y_e_spawn_3(3));
  Enemy_spawning_rngg_d13_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d13_n_0);
  Enemy_spawning_rngg_d14_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d14_n_0, CP => n_5, D => y_e_spawn_3(3), Q => y_e_spawn_1(1));
  Enemy_spawning_rngg_d14_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d14_n_0);
  Enemy_spawning_rngg_d15_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d15_n_0, CP => n_5, D => y_e_spawn_1(1), Q => y_e_spawn_3(1));
  Enemy_spawning_rngg_d15_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d15_n_0);
  Enemy_spawning_rngg_d16_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d16_n_0, CP => n_5, D => y_e_spawn_3(1), Q => y_e_spawn_1(0));
  Enemy_spawning_rngg_d16_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d16_n_0);
  Enemy_spawning_rngg_d1_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d1_n_0, CP => n_5, D => Enemy_spawning_rngg_xor_input, Q => y_e_spawn_5(8));
  Enemy_spawning_rngg_d1_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d1_n_0);
  Enemy_spawning_rngg_d2_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d2_n_0, CP => n_5, D => y_e_spawn_5(8), Q => y_e_spawn_1(8));
  Enemy_spawning_rngg_d2_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d2_n_0);
  Enemy_spawning_rngg_d3_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d3_n_0, CP => n_5, D => y_e_spawn_1(8), Q => y_e_spawn_2(7));
  Enemy_spawning_rngg_d3_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d3_n_0);
  Enemy_spawning_rngg_d4_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d4_n_0, CP => n_5, D => y_e_spawn_2(7), Q => y_e_spawn_1(7));
  Enemy_spawning_rngg_d4_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d4_n_0);
  Enemy_spawning_rngg_d5_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d5_n_0, CP => n_5, D => y_e_spawn_1(7), Q => y_e_spawn_4(7));
  Enemy_spawning_rngg_d5_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d5_n_0);
  Enemy_spawning_rngg_d6_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d6_n_0, CP => n_5, D => y_e_spawn_4(7), Q => y_e_spawn_1(5));
  Enemy_spawning_rngg_d6_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d6_n_0);
  Enemy_spawning_rngg_d7_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d7_n_0, CP => n_5, D => y_e_spawn_1(5), Q => y_e_spawn_3(7));
  Enemy_spawning_rngg_d7_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d7_n_0);
  Enemy_spawning_rngg_d8_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d8_n_0, CP => n_5, D => y_e_spawn_3(7), Q => y_e_spawn_1(4));
  Enemy_spawning_rngg_d8_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d8_n_0);
  Enemy_spawning_rngg_d9_q_reg : DFCNQD1BWP7T port map(CDN => Enemy_spawning_rngg_d9_n_0, CP => n_5, D => y_e_spawn_1(4), Q => y_e_spawn_2(3));
  Enemy_spawning_rngg_d9_g4 : INVD0BWP7T port map(I => reset, ZN => Enemy_spawning_rngg_d9_n_0);
  VGA_l044_count_reg_4 : DFCNQD1BWP7T port map(CDN => VGA_l044_n_0, CP => clk, D => VGA_l044_n_12, Q => VGA_draw_count4(4));
  VGA_l044_g82 : INR2D0BWP7T port map(A1 => VGA_enable4, B1 => VGA_l044_n_11, ZN => VGA_l044_n_12);
  VGA_l044_count_reg_3 : DFCNQD1BWP7T port map(CDN => VGA_l044_n_0, CP => clk, D => VGA_l044_n_10, Q => VGA_draw_count4(3));
  VGA_l044_g84 : MAOI22D0BWP7T port map(A1 => VGA_l044_n_8, A2 => VGA_draw_count4(4), B1 => VGA_l044_n_8, B2 => VGA_draw_count4(4), ZN => VGA_l044_n_11);
  VGA_l044_g85 : INR2D0BWP7T port map(A1 => VGA_enable4, B1 => VGA_l044_n_9, ZN => VGA_l044_n_10);
  VGA_l044_count_reg_2 : DFCNQD1BWP7T port map(CDN => VGA_l044_n_0, CP => clk, D => VGA_l044_n_7, Q => VGA_draw_count4(2));
  VGA_l044_g87 : MAOI22D0BWP7T port map(A1 => VGA_l044_n_4, A2 => VGA_draw_count4(3), B1 => VGA_l044_n_4, B2 => VGA_draw_count4(3), ZN => VGA_l044_n_9);
  VGA_l044_g88 : IND2D0BWP7T port map(A1 => VGA_l044_n_4, B1 => VGA_draw_count4(3), ZN => VGA_l044_n_8);
  VGA_l044_g89 : INR2D0BWP7T port map(A1 => VGA_enable4, B1 => VGA_l044_n_6, ZN => VGA_l044_n_7);
  VGA_l044_count_reg_1 : DFCNQD1BWP7T port map(CDN => VGA_l044_n_0, CP => clk, D => VGA_l044_n_5, Q => VGA_draw_count4(1));
  VGA_l044_g91 : MAOI22D0BWP7T port map(A1 => VGA_l044_n_1, A2 => VGA_draw_count4(2), B1 => VGA_l044_n_1, B2 => VGA_draw_count4(2), ZN => VGA_l044_n_6);
  VGA_l044_g92 : INR2D0BWP7T port map(A1 => VGA_enable4, B1 => VGA_l044_n_3, ZN => VGA_l044_n_5);
  VGA_l044_g93 : IND2D0BWP7T port map(A1 => VGA_l044_n_1, B1 => VGA_draw_count4(2), ZN => VGA_l044_n_4);
  VGA_l044_count_reg_0 : DFCNQD1BWP7T port map(CDN => VGA_l044_n_0, CP => clk, D => VGA_l044_n_2, Q => VGA_draw_count4(0));
  VGA_l044_g95 : XNR2D1BWP7T port map(A1 => VGA_draw_count4(0), A2 => VGA_draw_count4(1), ZN => VGA_l044_n_3);
  VGA_l044_g96 : INR2D0BWP7T port map(A1 => VGA_enable4, B1 => VGA_draw_count4(0), ZN => VGA_l044_n_2);
  VGA_l044_g97 : ND2D0BWP7T port map(A1 => VGA_draw_count4(0), A2 => VGA_draw_count4(1), ZN => VGA_l044_n_1);
  VGA_l044_g98 : INVD0BWP7T port map(I => reset, ZN => VGA_l044_n_0);
  VGA_l045_count_reg_4 : DFCNQD1BWP7T port map(CDN => VGA_l045_n_0, CP => clk, D => VGA_l045_n_12, Q => VGA_draw_count5(4));
  VGA_l045_g82 : INR2D0BWP7T port map(A1 => VGA_enable5, B1 => VGA_l045_n_11, ZN => VGA_l045_n_12);
  VGA_l045_count_reg_3 : DFCNQD1BWP7T port map(CDN => VGA_l045_n_0, CP => clk, D => VGA_l045_n_10, Q => VGA_draw_count5(3));
  VGA_l045_g84 : MAOI22D0BWP7T port map(A1 => VGA_l045_n_8, A2 => VGA_draw_count5(4), B1 => VGA_l045_n_8, B2 => VGA_draw_count5(4), ZN => VGA_l045_n_11);
  VGA_l045_g85 : INR2D0BWP7T port map(A1 => VGA_enable5, B1 => VGA_l045_n_9, ZN => VGA_l045_n_10);
  VGA_l045_count_reg_2 : DFCNQD1BWP7T port map(CDN => VGA_l045_n_0, CP => clk, D => VGA_l045_n_7, Q => VGA_draw_count5(2));
  VGA_l045_g87 : MAOI22D0BWP7T port map(A1 => VGA_l045_n_4, A2 => VGA_draw_count5(3), B1 => VGA_l045_n_4, B2 => VGA_draw_count5(3), ZN => VGA_l045_n_9);
  VGA_l045_g88 : IND2D0BWP7T port map(A1 => VGA_l045_n_4, B1 => VGA_draw_count5(3), ZN => VGA_l045_n_8);
  VGA_l045_g89 : INR2D0BWP7T port map(A1 => VGA_enable5, B1 => VGA_l045_n_6, ZN => VGA_l045_n_7);
  VGA_l045_count_reg_1 : DFCNQD1BWP7T port map(CDN => VGA_l045_n_0, CP => clk, D => VGA_l045_n_5, Q => VGA_draw_count5(1));
  VGA_l045_g91 : MAOI22D0BWP7T port map(A1 => VGA_l045_n_1, A2 => VGA_draw_count5(2), B1 => VGA_l045_n_1, B2 => VGA_draw_count5(2), ZN => VGA_l045_n_6);
  VGA_l045_g92 : INR2D0BWP7T port map(A1 => VGA_enable5, B1 => VGA_l045_n_3, ZN => VGA_l045_n_5);
  VGA_l045_g93 : IND2D0BWP7T port map(A1 => VGA_l045_n_1, B1 => VGA_draw_count5(2), ZN => VGA_l045_n_4);
  VGA_l045_count_reg_0 : DFCNQD1BWP7T port map(CDN => VGA_l045_n_0, CP => clk, D => VGA_l045_n_2, Q => VGA_draw_count5(0));
  VGA_l045_g95 : XNR2D1BWP7T port map(A1 => VGA_draw_count5(0), A2 => VGA_draw_count5(1), ZN => VGA_l045_n_3);
  VGA_l045_g96 : INR2D0BWP7T port map(A1 => VGA_enable5, B1 => VGA_draw_count5(0), ZN => VGA_l045_n_2);
  VGA_l045_g97 : ND2D0BWP7T port map(A1 => VGA_draw_count5(0), A2 => VGA_draw_count5(1), ZN => VGA_l045_n_1);
  VGA_l045_g98 : INVD0BWP7T port map(I => reset, ZN => VGA_l045_n_0);
  VGA_l046_count_reg_4 : DFCNQD1BWP7T port map(CDN => VGA_l046_n_0, CP => clk, D => VGA_l046_n_12, Q => VGA_draw_count6(4));
  VGA_l046_g82 : INR2D0BWP7T port map(A1 => VGA_enable6, B1 => VGA_l046_n_11, ZN => VGA_l046_n_12);
  VGA_l046_count_reg_3 : DFCNQD1BWP7T port map(CDN => VGA_l046_n_0, CP => clk, D => VGA_l046_n_10, Q => VGA_draw_count6(3));
  VGA_l046_g84 : MAOI22D0BWP7T port map(A1 => VGA_l046_n_8, A2 => VGA_draw_count6(4), B1 => VGA_l046_n_8, B2 => VGA_draw_count6(4), ZN => VGA_l046_n_11);
  VGA_l046_g85 : INR2D0BWP7T port map(A1 => VGA_enable6, B1 => VGA_l046_n_9, ZN => VGA_l046_n_10);
  VGA_l046_count_reg_2 : DFCNQD1BWP7T port map(CDN => VGA_l046_n_0, CP => clk, D => VGA_l046_n_7, Q => VGA_draw_count6(2));
  VGA_l046_g87 : MAOI22D0BWP7T port map(A1 => VGA_l046_n_4, A2 => VGA_draw_count6(3), B1 => VGA_l046_n_4, B2 => VGA_draw_count6(3), ZN => VGA_l046_n_9);
  VGA_l046_g88 : IND2D0BWP7T port map(A1 => VGA_l046_n_4, B1 => VGA_draw_count6(3), ZN => VGA_l046_n_8);
  VGA_l046_g89 : INR2D0BWP7T port map(A1 => VGA_enable6, B1 => VGA_l046_n_6, ZN => VGA_l046_n_7);
  VGA_l046_count_reg_1 : DFCNQD1BWP7T port map(CDN => VGA_l046_n_0, CP => clk, D => VGA_l046_n_5, Q => VGA_draw_count6(1));
  VGA_l046_g91 : MAOI22D0BWP7T port map(A1 => VGA_l046_n_1, A2 => VGA_draw_count6(2), B1 => VGA_l046_n_1, B2 => VGA_draw_count6(2), ZN => VGA_l046_n_6);
  VGA_l046_g92 : INR2D0BWP7T port map(A1 => VGA_enable6, B1 => VGA_l046_n_3, ZN => VGA_l046_n_5);
  VGA_l046_g93 : IND2D0BWP7T port map(A1 => VGA_l046_n_1, B1 => VGA_draw_count6(2), ZN => VGA_l046_n_4);
  VGA_l046_count_reg_0 : DFCNQD1BWP7T port map(CDN => VGA_l046_n_0, CP => clk, D => VGA_l046_n_2, Q => VGA_draw_count6(0));
  VGA_l046_g95 : XNR2D1BWP7T port map(A1 => VGA_draw_count6(0), A2 => VGA_draw_count6(1), ZN => VGA_l046_n_3);
  VGA_l046_g96 : INR2D0BWP7T port map(A1 => VGA_enable6, B1 => VGA_draw_count6(0), ZN => VGA_l046_n_2);
  VGA_l046_g97 : ND2D0BWP7T port map(A1 => VGA_draw_count6(0), A2 => VGA_draw_count6(1), ZN => VGA_l046_n_1);
  VGA_l046_g98 : INVD0BWP7T port map(I => reset, ZN => VGA_l046_n_0);
  Enemy_spawning_en51_decider_reg : DFQD1BWP7T port map(CP => clk, D => Enemy_spawning_en51_n_3, Q => spawn_or_not_e5);
  Enemy_spawning_en51_g143 : NR4D0BWP7T port map(A1 => Enemy_spawning_en51_n_2, A2 => Enemy_spawning_en51_n_1, A3 => Enemy_spawning_en51_n_0, A4 => e_5, ZN => Enemy_spawning_en51_n_3);
  Enemy_spawning_en51_g144 : ND4D0BWP7T port map(A1 => y_e_spawn_2(3), A2 => y_e_spawn_1(4), A3 => y_e_spawn_1(8), A4 => y_e_spawn_5(8), ZN => Enemy_spawning_en51_n_2);
  Enemy_spawning_en51_g145 : ND2D0BWP7T port map(A1 => y_e_spawn_1(5), A2 => y_e_spawn_3(7), ZN => Enemy_spawning_en51_n_1);
  Enemy_spawning_en51_g146 : ND2D0BWP7T port map(A1 => y_e_spawn_1(1), A2 => n_5, ZN => Enemy_spawning_en51_n_0);
  VGA_l047_count_reg_4 : DFCNQD1BWP7T port map(CDN => VGA_l047_n_0, CP => clk, D => VGA_l047_n_12, Q => VGA_draw_count7(4));
  VGA_l047_g82 : INR2D0BWP7T port map(A1 => VGA_enable7, B1 => VGA_l047_n_11, ZN => VGA_l047_n_12);
  VGA_l047_count_reg_3 : DFCNQD1BWP7T port map(CDN => VGA_l047_n_0, CP => clk, D => VGA_l047_n_10, Q => VGA_draw_count7(3));
  VGA_l047_g84 : MAOI22D0BWP7T port map(A1 => VGA_l047_n_8, A2 => VGA_draw_count7(4), B1 => VGA_l047_n_8, B2 => VGA_draw_count7(4), ZN => VGA_l047_n_11);
  VGA_l047_g85 : INR2D0BWP7T port map(A1 => VGA_enable7, B1 => VGA_l047_n_9, ZN => VGA_l047_n_10);
  VGA_l047_count_reg_2 : DFCNQD1BWP7T port map(CDN => VGA_l047_n_0, CP => clk, D => VGA_l047_n_7, Q => VGA_draw_count7(2));
  VGA_l047_g87 : MAOI22D0BWP7T port map(A1 => VGA_l047_n_4, A2 => VGA_draw_count7(3), B1 => VGA_l047_n_4, B2 => VGA_draw_count7(3), ZN => VGA_l047_n_9);
  VGA_l047_g88 : IND2D0BWP7T port map(A1 => VGA_l047_n_4, B1 => VGA_draw_count7(3), ZN => VGA_l047_n_8);
  VGA_l047_g89 : INR2D0BWP7T port map(A1 => VGA_enable7, B1 => VGA_l047_n_6, ZN => VGA_l047_n_7);
  VGA_l047_count_reg_1 : DFCNQD1BWP7T port map(CDN => VGA_l047_n_0, CP => clk, D => VGA_l047_n_5, Q => VGA_draw_count7(1));
  VGA_l047_g91 : MAOI22D0BWP7T port map(A1 => VGA_l047_n_1, A2 => VGA_draw_count7(2), B1 => VGA_l047_n_1, B2 => VGA_draw_count7(2), ZN => VGA_l047_n_6);
  VGA_l047_g92 : INR2D0BWP7T port map(A1 => VGA_enable7, B1 => VGA_l047_n_3, ZN => VGA_l047_n_5);
  VGA_l047_g93 : IND2D0BWP7T port map(A1 => VGA_l047_n_1, B1 => VGA_draw_count7(2), ZN => VGA_l047_n_4);
  VGA_l047_count_reg_0 : DFCNQD1BWP7T port map(CDN => VGA_l047_n_0, CP => clk, D => VGA_l047_n_2, Q => VGA_draw_count7(0));
  VGA_l047_g95 : XNR2D1BWP7T port map(A1 => VGA_draw_count7(0), A2 => VGA_draw_count7(1), ZN => VGA_l047_n_3);
  VGA_l047_g96 : INR2D0BWP7T port map(A1 => VGA_enable7, B1 => VGA_draw_count7(0), ZN => VGA_l047_n_2);
  VGA_l047_g97 : ND2D0BWP7T port map(A1 => VGA_draw_count7(0), A2 => VGA_draw_count7(1), ZN => VGA_l047_n_1);
  VGA_l047_g98 : INVD0BWP7T port map(I => reset, ZN => VGA_l047_n_0);
  VGA_l048_count_reg_4 : DFCNQD1BWP7T port map(CDN => VGA_l048_n_0, CP => clk, D => VGA_l048_n_12, Q => VGA_draw_count8(4));
  VGA_l048_g82 : INR2D0BWP7T port map(A1 => VGA_enable8, B1 => VGA_l048_n_11, ZN => VGA_l048_n_12);
  VGA_l048_count_reg_3 : DFCNQD1BWP7T port map(CDN => VGA_l048_n_0, CP => clk, D => VGA_l048_n_10, Q => VGA_draw_count8(3));
  VGA_l048_g84 : MAOI22D0BWP7T port map(A1 => VGA_l048_n_8, A2 => VGA_draw_count8(4), B1 => VGA_l048_n_8, B2 => VGA_draw_count8(4), ZN => VGA_l048_n_11);
  VGA_l048_g85 : INR2D0BWP7T port map(A1 => VGA_enable8, B1 => VGA_l048_n_9, ZN => VGA_l048_n_10);
  VGA_l048_count_reg_2 : DFCNQD1BWP7T port map(CDN => VGA_l048_n_0, CP => clk, D => VGA_l048_n_7, Q => VGA_draw_count8(2));
  VGA_l048_g87 : MAOI22D0BWP7T port map(A1 => VGA_l048_n_4, A2 => VGA_draw_count8(3), B1 => VGA_l048_n_4, B2 => VGA_draw_count8(3), ZN => VGA_l048_n_9);
  VGA_l048_g88 : IND2D0BWP7T port map(A1 => VGA_l048_n_4, B1 => VGA_draw_count8(3), ZN => VGA_l048_n_8);
  VGA_l048_g89 : INR2D0BWP7T port map(A1 => VGA_enable8, B1 => VGA_l048_n_6, ZN => VGA_l048_n_7);
  VGA_l048_count_reg_1 : DFCNQD1BWP7T port map(CDN => VGA_l048_n_0, CP => clk, D => VGA_l048_n_5, Q => VGA_draw_count8(1));
  VGA_l048_g91 : MAOI22D0BWP7T port map(A1 => VGA_l048_n_1, A2 => VGA_draw_count8(2), B1 => VGA_l048_n_1, B2 => VGA_draw_count8(2), ZN => VGA_l048_n_6);
  VGA_l048_g92 : INR2D0BWP7T port map(A1 => VGA_enable8, B1 => VGA_l048_n_3, ZN => VGA_l048_n_5);
  VGA_l048_g93 : IND2D0BWP7T port map(A1 => VGA_l048_n_1, B1 => VGA_draw_count8(2), ZN => VGA_l048_n_4);
  VGA_l048_count_reg_0 : DFCNQD1BWP7T port map(CDN => VGA_l048_n_0, CP => clk, D => VGA_l048_n_2, Q => VGA_draw_count8(0));
  VGA_l048_g95 : XNR2D1BWP7T port map(A1 => VGA_draw_count8(0), A2 => VGA_draw_count8(1), ZN => VGA_l048_n_3);
  VGA_l048_g96 : INR2D0BWP7T port map(A1 => VGA_enable8, B1 => VGA_draw_count8(0), ZN => VGA_l048_n_2);
  VGA_l048_g97 : ND2D0BWP7T port map(A1 => VGA_draw_count8(0), A2 => VGA_draw_count8(1), ZN => VGA_l048_n_1);
  VGA_l048_g98 : INVD0BWP7T port map(I => reset, ZN => VGA_l048_n_0);
  VGA_l0410_count_reg_4 : DFCNQD1BWP7T port map(CDN => VGA_l0410_n_0, CP => clk, D => VGA_l0410_n_12, Q => VGA_draw_count10(4));
  VGA_l0410_g82 : INR2D0BWP7T port map(A1 => VGA_enable10, B1 => VGA_l0410_n_11, ZN => VGA_l0410_n_12);
  VGA_l0410_count_reg_3 : DFCNQD1BWP7T port map(CDN => VGA_l0410_n_0, CP => clk, D => VGA_l0410_n_10, Q => VGA_draw_count10(3));
  VGA_l0410_g84 : MAOI22D0BWP7T port map(A1 => VGA_l0410_n_8, A2 => VGA_draw_count10(4), B1 => VGA_l0410_n_8, B2 => VGA_draw_count10(4), ZN => VGA_l0410_n_11);
  VGA_l0410_g85 : INR2D0BWP7T port map(A1 => VGA_enable10, B1 => VGA_l0410_n_9, ZN => VGA_l0410_n_10);
  VGA_l0410_count_reg_2 : DFCNQD1BWP7T port map(CDN => VGA_l0410_n_0, CP => clk, D => VGA_l0410_n_7, Q => VGA_draw_count10(2));
  VGA_l0410_g87 : MAOI22D0BWP7T port map(A1 => VGA_l0410_n_4, A2 => VGA_draw_count10(3), B1 => VGA_l0410_n_4, B2 => VGA_draw_count10(3), ZN => VGA_l0410_n_9);
  VGA_l0410_g88 : IND2D0BWP7T port map(A1 => VGA_l0410_n_4, B1 => VGA_draw_count10(3), ZN => VGA_l0410_n_8);
  VGA_l0410_g89 : INR2D0BWP7T port map(A1 => VGA_enable10, B1 => VGA_l0410_n_6, ZN => VGA_l0410_n_7);
  VGA_l0410_count_reg_1 : DFCNQD1BWP7T port map(CDN => VGA_l0410_n_0, CP => clk, D => VGA_l0410_n_5, Q => VGA_draw_count10(1));
  VGA_l0410_g91 : MAOI22D0BWP7T port map(A1 => VGA_l0410_n_1, A2 => VGA_draw_count10(2), B1 => VGA_l0410_n_1, B2 => VGA_draw_count10(2), ZN => VGA_l0410_n_6);
  VGA_l0410_g92 : INR2D0BWP7T port map(A1 => VGA_enable10, B1 => VGA_l0410_n_3, ZN => VGA_l0410_n_5);
  VGA_l0410_g93 : IND2D0BWP7T port map(A1 => VGA_l0410_n_1, B1 => VGA_draw_count10(2), ZN => VGA_l0410_n_4);
  VGA_l0410_count_reg_0 : DFCNQD1BWP7T port map(CDN => VGA_l0410_n_0, CP => clk, D => VGA_l0410_n_2, Q => VGA_draw_count10(0));
  VGA_l0410_g95 : XNR2D1BWP7T port map(A1 => VGA_draw_count10(0), A2 => VGA_draw_count10(1), ZN => VGA_l0410_n_3);
  VGA_l0410_g96 : INR2D0BWP7T port map(A1 => VGA_enable10, B1 => VGA_draw_count10(0), ZN => VGA_l0410_n_2);
  VGA_l0410_g97 : ND2D0BWP7T port map(A1 => VGA_draw_count10(0), A2 => VGA_draw_count10(1), ZN => VGA_l0410_n_1);
  VGA_l0410_g98 : INVD0BWP7T port map(I => reset, ZN => VGA_l0410_n_0);
  VGA_l049_count_reg_4 : DFCNQD1BWP7T port map(CDN => VGA_l049_n_0, CP => clk, D => VGA_l049_n_12, Q => VGA_draw_count9(4));
  VGA_l049_g82 : INR2D0BWP7T port map(A1 => VGA_enable9, B1 => VGA_l049_n_11, ZN => VGA_l049_n_12);
  VGA_l049_count_reg_3 : DFCNQD1BWP7T port map(CDN => VGA_l049_n_0, CP => clk, D => VGA_l049_n_10, Q => VGA_draw_count9(3));
  VGA_l049_g84 : MAOI22D0BWP7T port map(A1 => VGA_l049_n_8, A2 => VGA_draw_count9(4), B1 => VGA_l049_n_8, B2 => VGA_draw_count9(4), ZN => VGA_l049_n_11);
  VGA_l049_g85 : INR2D0BWP7T port map(A1 => VGA_enable9, B1 => VGA_l049_n_9, ZN => VGA_l049_n_10);
  VGA_l049_count_reg_2 : DFCNQD1BWP7T port map(CDN => VGA_l049_n_0, CP => clk, D => VGA_l049_n_7, Q => VGA_draw_count9(2));
  VGA_l049_g87 : MAOI22D0BWP7T port map(A1 => VGA_l049_n_4, A2 => VGA_draw_count9(3), B1 => VGA_l049_n_4, B2 => VGA_draw_count9(3), ZN => VGA_l049_n_9);
  VGA_l049_g88 : IND2D0BWP7T port map(A1 => VGA_l049_n_4, B1 => VGA_draw_count9(3), ZN => VGA_l049_n_8);
  VGA_l049_g89 : INR2D0BWP7T port map(A1 => VGA_enable9, B1 => VGA_l049_n_6, ZN => VGA_l049_n_7);
  VGA_l049_count_reg_1 : DFCNQD1BWP7T port map(CDN => VGA_l049_n_0, CP => clk, D => VGA_l049_n_5, Q => VGA_draw_count9(1));
  VGA_l049_g91 : MAOI22D0BWP7T port map(A1 => VGA_l049_n_1, A2 => VGA_draw_count9(2), B1 => VGA_l049_n_1, B2 => VGA_draw_count9(2), ZN => VGA_l049_n_6);
  VGA_l049_g92 : INR2D0BWP7T port map(A1 => VGA_enable9, B1 => VGA_l049_n_3, ZN => VGA_l049_n_5);
  VGA_l049_g93 : IND2D0BWP7T port map(A1 => VGA_l049_n_1, B1 => VGA_draw_count9(2), ZN => VGA_l049_n_4);
  VGA_l049_count_reg_0 : DFCNQD1BWP7T port map(CDN => VGA_l049_n_0, CP => clk, D => VGA_l049_n_2, Q => VGA_draw_count9(0));
  VGA_l049_g95 : XNR2D1BWP7T port map(A1 => VGA_draw_count9(0), A2 => VGA_draw_count9(1), ZN => VGA_l049_n_3);
  VGA_l049_g96 : INR2D0BWP7T port map(A1 => VGA_enable9, B1 => VGA_draw_count9(0), ZN => VGA_l049_n_2);
  VGA_l049_g97 : ND2D0BWP7T port map(A1 => VGA_draw_count9(0), A2 => VGA_draw_count9(1), ZN => VGA_l049_n_1);
  VGA_l049_g98 : INVD0BWP7T port map(I => reset, ZN => VGA_l049_n_0);
  VGA_l051_g2479 : AO31D0BWP7T port map(A1 => VGA_l051_n_77, A2 => VGA_l051_n_76, A3 => VGA_draw_count1(0), B => VGA_b1, Z => VGA_g1);
  VGA_l051_g2480 : OA21D0BWP7T port map(A1 => VGA_l051_n_79, A2 => VGA_l051_n_39, B => VGA_enable1, Z => VGA_r1);
  VGA_l051_g2481 : AO32D0BWP7T port map(A1 => VGA_l051_n_77, A2 => VGA_l051_n_76, A3 => VGA_l051_n_17, B1 => VGA_l051_n_78, B2 => VGA_l051_n_39, Z => VGA_b1);
  VGA_l051_g2482 : IND2D0BWP7T port map(A1 => VGA_l051_n_77, B1 => VGA_l051_n_75, ZN => VGA_enable1);
  VGA_l051_g2483 : MOAI22D0BWP7T port map(A1 => VGA_l051_n_4, A2 => VGA_draw_count1(2), B1 => VGA_l051_n_76, B2 => VGA_l051_n_73, ZN => VGA_l051_n_79);
  VGA_l051_g2484 : ND2D0BWP7T port map(A1 => VGA_l051_n_76, A2 => VGA_l051_n_75, ZN => VGA_l051_n_78);
  VGA_l051_g2485 : IAO21D0BWP7T port map(A1 => VGA_l051_n_74, A2 => VGA_l051_n_0, B => VGA_l051_n_72, ZN => VGA_l051_n_77);
  VGA_l051_g2486 : IND2D0BWP7T port map(A1 => VGA_l051_n_72, B1 => VGA_l051_n_74, ZN => VGA_l051_n_76);
  VGA_l051_g2487 : OR2D0BWP7T port map(A1 => VGA_l051_n_73, A2 => VGA_l051_n_72, Z => VGA_l051_n_75);
  VGA_l051_g2489 : NR4D0BWP7T port map(A1 => VGA_l051_n_71, A2 => VGA_l051_n_47, A3 => VGA_l051_n_29, A4 => VGA_l051_n_27, ZN => VGA_l051_n_74);
  VGA_l051_g2490 : ND4D0BWP7T port map(A1 => VGA_l051_n_70, A2 => VGA_l051_n_35, A3 => VGA_l051_n_27, A4 => VGA_l051_n_25, ZN => VGA_l051_n_73);
  VGA_l051_g2491 : ND4D0BWP7T port map(A1 => VGA_l051_n_67, A2 => VGA_l051_n_69, A3 => VGA_l051_n_55, A4 => VGA_l051_n_49, ZN => VGA_l051_n_72);
  VGA_l051_g2492 : OAI211D0BWP7T port map(A1 => VGA_l051_n_12, A2 => VGA_l051_n_30, B => VGA_l051_n_68, C => VGA_l051_n_56, ZN => VGA_l051_n_71);
  VGA_l051_g2493 : NR4D0BWP7T port map(A1 => VGA_l051_n_64, A2 => VGA_l051_n_57, A3 => VGA_l051_n_28, A4 => VGA_l051_n_29, ZN => VGA_l051_n_70);
  VGA_l051_g2494 : AOI211D0BWP7T port map(A1 => VGA_l051_n_7, A2 => VGA_l051_n_10, B => VGA_l051_n_66, C => VGA_l051_n_51, ZN => VGA_l051_n_69);
  VGA_l051_g2495 : NR4D0BWP7T port map(A1 => VGA_l051_n_61, A2 => VGA_l051_n_63, A3 => VGA_l051_n_53, A4 => VGA_l051_n_57, ZN => VGA_l051_n_68);
  VGA_l051_g2496 : OAI31D0BWP7T port map(A1 => VGA_l051_n_15, A2 => VGA_l051_n_34, A3 => VGA_l051_n_60, B => VGA_l051_n_65, ZN => VGA_l051_n_67);
  VGA_l051_g2497 : AOI22D0BWP7T port map(A1 => VGA_l051_n_62, A2 => VGA_l051_n_50, B1 => VGA_l051_n_33, B2 => VGA_l051_n_9, ZN => VGA_l051_n_66);
  VGA_l051_g2498 : OA32D0BWP7T port map(A1 => VGA_l051_n_20, A2 => VGA_l051_n_33, A3 => VGA_l051_n_1, B1 => VGA_l051_n_60, B2 => VGA_l051_n_58, Z => VGA_l051_n_65);
  VGA_l051_g2499 : OR3D0BWP7T port map(A1 => VGA_l051_n_30, A2 => VGA_l051_n_52, A3 => VGA_l051_n_63, Z => VGA_l051_n_64);
  VGA_l051_g2500 : OAI211D0BWP7T port map(A1 => VGA_l051_n_5, A2 => VGA_l051_n_11, B => VGA_l051_n_45, C => VGA_l051_n_19, ZN => VGA_l051_n_62);
  VGA_l051_g2501 : OAI221D0BWP7T port map(A1 => VGA_l051_n_35, A2 => VGA_l051_n_22, B1 => VGA_l051_n_16, B2 => VGA_l051_n_26, C => VGA_l051_n_48, ZN => VGA_l051_n_61);
  VGA_l051_g2502 : OAI211D0BWP7T port map(A1 => VGA_l051_n_18, A2 => VGA_l051_n_38, B => VGA_l051_n_46, C => VGA_l051_n_54, ZN => VGA_l051_n_63);
  VGA_l051_g2503 : MOAI22D0BWP7T port map(A1 => VGA_l051_n_25, A2 => y_pos_b1(1), B1 => VGA_l051_n_47, B2 => y_pos_b1(1), ZN => VGA_l051_n_59);
  VGA_l051_g2504 : OAI211D0BWP7T port map(A1 => VGA_l051_n_11, A2 => VGA_l051_n_36, B => VGA_l051_n_43, C => VGA_l051_n_44, ZN => VGA_l051_n_58);
  VGA_l051_g2505 : AO21D0BWP7T port map(A1 => VGA_l051_n_33, A2 => VGA_l051_n_20, B => VGA_l051_n_1, Z => VGA_l051_n_60);
  VGA_l051_g2506 : AOI22D0BWP7T port map(A1 => VGA_l051_n_30, A2 => VGA_l051_n_12, B1 => VGA_l051_n_41, B2 => VGA_y(1), ZN => VGA_l051_n_56);
  VGA_l051_g2507 : AOI22D0BWP7T port map(A1 => VGA_l051_n_37, A2 => VGA_l051_n_13, B1 => VGA_l051_n_2, B2 => x_pos_b1(8), ZN => VGA_l051_n_55);
  VGA_l051_g2508 : MAOI22D0BWP7T port map(A1 => VGA_l051_n_21, A2 => VGA_y(9), B1 => VGA_l051_n_21, B2 => VGA_y(9), ZN => VGA_l051_n_54);
  VGA_l051_g2509 : MOAI22D0BWP7T port map(A1 => VGA_l051_n_28, A2 => VGA_l051_n_14, B1 => VGA_l051_n_28, B2 => VGA_l051_n_14, ZN => VGA_l051_n_53);
  VGA_l051_g2510 : MAOI22D0BWP7T port map(A1 => VGA_l051_n_31, A2 => VGA_l051_n_23, B1 => VGA_l051_n_31, B2 => VGA_l051_n_23, ZN => VGA_l051_n_57);
  VGA_l051_g2511 : MOAI22D0BWP7T port map(A1 => VGA_l051_n_26, A2 => VGA_y(5), B1 => VGA_l051_n_26, B2 => VGA_y(5), ZN => VGA_l051_n_52);
  VGA_l051_g2512 : OAI22D0BWP7T port map(A1 => VGA_l051_n_40, A2 => VGA_l051_n_6, B1 => VGA_l051_n_32, B2 => VGA_l051_n_8, ZN => VGA_l051_n_51);
  VGA_l051_g2513 : MAOI22D0BWP7T port map(A1 => VGA_l051_n_34, A2 => VGA_l051_n_24, B1 => VGA_l051_n_33, B2 => VGA_l051_n_9, ZN => VGA_l051_n_50);
  VGA_l051_g2514 : MAOI22D0BWP7T port map(A1 => VGA_l051_n_32, A2 => VGA_l051_n_8, B1 => VGA_l051_n_7, B2 => VGA_l051_n_10, ZN => VGA_l051_n_49);
  VGA_l051_g2515 : AOI22D0BWP7T port map(A1 => VGA_l051_n_26, A2 => VGA_l051_n_16, B1 => VGA_l051_n_35, B2 => VGA_l051_n_22, ZN => VGA_l051_n_48);
  VGA_l051_g2517 : ND2D0BWP7T port map(A1 => VGA_l051_n_38, A2 => VGA_l051_n_18, ZN => VGA_l051_n_46);
  VGA_l051_g2518 : IND2D0BWP7T port map(A1 => VGA_l051_n_34, B1 => VGA_l051_n_15, ZN => VGA_l051_n_45);
  VGA_l051_g2519 : NR2D0BWP7T port map(A1 => VGA_l051_n_41, A2 => VGA_y(1), ZN => VGA_l051_n_47);
  VGA_l051_g2520 : ND2D0BWP7T port map(A1 => VGA_l051_n_34, A2 => VGA_l051_n_15, ZN => VGA_l051_n_44);
  VGA_l051_g2521 : AO21D0BWP7T port map(A1 => VGA_l051_n_36, A2 => VGA_l051_n_19, B => VGA_l051_n_5, Z => VGA_l051_n_43);
  VGA_l051_g2522 : CKXOR2D0BWP7T port map(A1 => VGA_y(0), A2 => VGA_l051_n_27, Z => VGA_l051_n_42);
  VGA_l051_g2525 : CKND1BWP7T port map(I => VGA_l051_n_25, ZN => VGA_l051_n_41);
  VGA_l051_g2526 : MOAI22D0BWP7T port map(A1 => VGA_x(6), A2 => x_pos_b1(6), B1 => VGA_x(6), B2 => x_pos_b1(6), ZN => VGA_l051_n_40);
  VGA_l051_g2527 : OA21D0BWP7T port map(A1 => VGA_l051_n_4, A2 => VGA_draw_count1(1), B => VGA_l051_n_17, Z => VGA_l051_n_39);
  VGA_l051_g2528 : MOAI22D0BWP7T port map(A1 => VGA_y(8), A2 => y_pos_b1(8), B1 => VGA_y(8), B2 => y_pos_b1(8), ZN => VGA_l051_n_38);
  VGA_l051_g2529 : MOAI22D0BWP7T port map(A1 => VGA_x(5), A2 => x_pos_b1(5), B1 => VGA_x(5), B2 => x_pos_b1(5), ZN => VGA_l051_n_37);
  VGA_l051_g2530 : AN2D1BWP7T port map(A1 => VGA_l051_n_15, A2 => VGA_l051_n_24, Z => VGA_l051_n_36);
  VGA_l051_g2531 : AO21D0BWP7T port map(A1 => VGA_l051_n_3, A2 => y_pos_b1(5), B => VGA_l051_n_16, Z => VGA_l051_n_35);
  VGA_l051_g2532 : MOAI22D0BWP7T port map(A1 => VGA_x(3), A2 => x_pos_b1(3), B1 => VGA_x(3), B2 => x_pos_b1(3), ZN => VGA_l051_n_34);
  VGA_l051_g2533 : MAOI22D0BWP7T port map(A1 => VGA_x(4), A2 => x_pos_b1(4), B1 => VGA_x(4), B2 => x_pos_b1(4), ZN => VGA_l051_n_33);
  VGA_l051_g2535 : MAOI22D0BWP7T port map(A1 => VGA_x(7), A2 => x_pos_b1(7), B1 => VGA_x(7), B2 => x_pos_b1(7), ZN => VGA_l051_n_32);
  VGA_l051_g2536 : MAOI22D0BWP7T port map(A1 => VGA_y(7), A2 => y_pos_b1(7), B1 => VGA_y(7), B2 => y_pos_b1(7), ZN => VGA_l051_n_31);
  VGA_l051_g2537 : MAOI22D0BWP7T port map(A1 => VGA_y(3), A2 => y_pos_b1(3), B1 => VGA_y(3), B2 => y_pos_b1(3), ZN => VGA_l051_n_30);
  VGA_l051_g2538 : MAOI22D0BWP7T port map(A1 => VGA_y(0), A2 => y_pos_b1(0), B1 => VGA_y(0), B2 => y_pos_b1(0), ZN => VGA_l051_n_29);
  VGA_l051_g2539 : MAOI22D0BWP7T port map(A1 => VGA_y(4), A2 => y_pos_b1(4), B1 => VGA_y(4), B2 => y_pos_b1(4), ZN => VGA_l051_n_28);
  VGA_l051_g2540 : MOAI22D0BWP7T port map(A1 => VGA_y(1), A2 => y_pos_b1(1), B1 => VGA_y(1), B2 => y_pos_b1(1), ZN => VGA_l051_n_27);
  VGA_l051_g2541 : MAOI22D0BWP7T port map(A1 => VGA_y(6), A2 => y_pos_b1(6), B1 => VGA_y(6), B2 => y_pos_b1(6), ZN => VGA_l051_n_26);
  VGA_l051_g2542 : MOAI22D0BWP7T port map(A1 => VGA_y(2), A2 => y_pos_b1(2), B1 => VGA_y(2), B2 => y_pos_b1(2), ZN => VGA_l051_n_25);
  VGA_l051_g2543 : IND2D0BWP7T port map(A1 => x_pos_b1(2), B1 => VGA_x(2), ZN => VGA_l051_n_24);
  VGA_l051_g2544 : INR2D0BWP7T port map(A1 => y_pos_b1(6), B1 => VGA_y(6), ZN => VGA_l051_n_23);
  VGA_l051_g2545 : INR2D0BWP7T port map(A1 => y_pos_b1(4), B1 => VGA_y(4), ZN => VGA_l051_n_22);
  VGA_l051_g2546 : IND2D0BWP7T port map(A1 => VGA_y(8), B1 => y_pos_b1(8), ZN => VGA_l051_n_21);
  VGA_l051_g2547 : INR2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_b1(3), ZN => VGA_l051_n_20);
  VGA_l051_g2548 : IND2D0BWP7T port map(A1 => x_pos_b1(1), B1 => VGA_x(1), ZN => VGA_l051_n_19);
  VGA_l051_g2549 : INR2D0BWP7T port map(A1 => y_pos_b1(7), B1 => VGA_y(7), ZN => VGA_l051_n_18);
  VGA_l051_g2550 : OR2D0BWP7T port map(A1 => VGA_draw_count1(2), A2 => VGA_draw_count1(1), Z => VGA_l051_n_17);
  VGA_l051_g2551 : NR2D0BWP7T port map(A1 => VGA_l051_n_3, A2 => y_pos_b1(5), ZN => VGA_l051_n_16);
  VGA_l051_g2552 : IND2D0BWP7T port map(A1 => VGA_x(2), B1 => x_pos_b1(2), ZN => VGA_l051_n_15);
  VGA_l051_g2553 : IND2D0BWP7T port map(A1 => VGA_y(3), B1 => y_pos_b1(3), ZN => VGA_l051_n_14);
  VGA_l051_g2554 : INR2D0BWP7T port map(A1 => x_pos_b1(4), B1 => VGA_x(4), ZN => VGA_l051_n_13);
  VGA_l051_g2555 : IND2D0BWP7T port map(A1 => VGA_y(2), B1 => y_pos_b1(2), ZN => VGA_l051_n_12);
  VGA_l051_g2556 : INR2D0BWP7T port map(A1 => x_pos_b1(1), B1 => VGA_x(1), ZN => VGA_l051_n_11);
  VGA_l051_g2557 : IND2D0BWP7T port map(A1 => x_pos_b1(8), B1 => VGA_x(8), ZN => VGA_l051_n_10);
  VGA_l051_g2558 : IND2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_b1(3), ZN => VGA_l051_n_9);
  VGA_l051_g2559 : INR2D0BWP7T port map(A1 => VGA_x(6), B1 => x_pos_b1(6), ZN => VGA_l051_n_8);
  VGA_l051_g2560 : INR2D0BWP7T port map(A1 => x_pos_b1(7), B1 => VGA_x(7), ZN => VGA_l051_n_7);
  VGA_l051_g2561 : IND2D0BWP7T port map(A1 => VGA_x(5), B1 => x_pos_b1(5), ZN => VGA_l051_n_6);
  VGA_l051_g2562 : IND2D0BWP7T port map(A1 => x_pos_b1(0), B1 => VGA_x(0), ZN => VGA_l051_n_5);
  VGA_l051_g2563 : CKND1BWP7T port map(I => VGA_draw_count1(0), ZN => VGA_l051_n_4);
  VGA_l051_g2564 : CKND1BWP7T port map(I => VGA_y(5), ZN => VGA_l051_n_3);
  VGA_l051_g2565 : CKND1BWP7T port map(I => VGA_x(8), ZN => VGA_l051_n_2);
  VGA_l051_g2 : MOAI22D0BWP7T port map(A1 => VGA_l051_n_37, A2 => VGA_l051_n_13, B1 => VGA_l051_n_40, B2 => VGA_l051_n_6, ZN => VGA_l051_n_1);
  VGA_l051_g2566 : INR4D0BWP7T port map(A1 => VGA_l051_n_29, B1 => VGA_l051_n_71, B2 => VGA_l051_n_59, B3 => VGA_l051_n_42, ZN => VGA_l051_n_0);
  VGA_l052_g2479 : AO31D0BWP7T port map(A1 => VGA_l052_n_77, A2 => VGA_l052_n_76, A3 => VGA_draw_count2(0), B => VGA_b2, Z => VGA_g2);
  VGA_l052_g2480 : OA21D0BWP7T port map(A1 => VGA_l052_n_79, A2 => VGA_l052_n_39, B => VGA_enable2, Z => VGA_r2);
  VGA_l052_g2481 : AO32D0BWP7T port map(A1 => VGA_l052_n_77, A2 => VGA_l052_n_76, A3 => VGA_l052_n_17, B1 => VGA_l052_n_78, B2 => VGA_l052_n_39, Z => VGA_b2);
  VGA_l052_g2482 : IND2D0BWP7T port map(A1 => VGA_l052_n_77, B1 => VGA_l052_n_75, ZN => VGA_enable2);
  VGA_l052_g2483 : MOAI22D0BWP7T port map(A1 => VGA_l052_n_4, A2 => VGA_draw_count2(2), B1 => VGA_l052_n_76, B2 => VGA_l052_n_73, ZN => VGA_l052_n_79);
  VGA_l052_g2484 : ND2D0BWP7T port map(A1 => VGA_l052_n_76, A2 => VGA_l052_n_75, ZN => VGA_l052_n_78);
  VGA_l052_g2485 : IAO21D0BWP7T port map(A1 => VGA_l052_n_74, A2 => VGA_l052_n_0, B => VGA_l052_n_72, ZN => VGA_l052_n_77);
  VGA_l052_g2486 : IND2D0BWP7T port map(A1 => VGA_l052_n_72, B1 => VGA_l052_n_74, ZN => VGA_l052_n_76);
  VGA_l052_g2487 : OR2D0BWP7T port map(A1 => VGA_l052_n_73, A2 => VGA_l052_n_72, Z => VGA_l052_n_75);
  VGA_l052_g2489 : NR4D0BWP7T port map(A1 => VGA_l052_n_71, A2 => VGA_l052_n_47, A3 => VGA_l052_n_29, A4 => VGA_l052_n_27, ZN => VGA_l052_n_74);
  VGA_l052_g2490 : ND4D0BWP7T port map(A1 => VGA_l052_n_70, A2 => VGA_l052_n_35, A3 => VGA_l052_n_27, A4 => VGA_l052_n_25, ZN => VGA_l052_n_73);
  VGA_l052_g2491 : ND4D0BWP7T port map(A1 => VGA_l052_n_67, A2 => VGA_l052_n_69, A3 => VGA_l052_n_55, A4 => VGA_l052_n_49, ZN => VGA_l052_n_72);
  VGA_l052_g2492 : OAI211D0BWP7T port map(A1 => VGA_l052_n_12, A2 => VGA_l052_n_30, B => VGA_l052_n_68, C => VGA_l052_n_56, ZN => VGA_l052_n_71);
  VGA_l052_g2493 : NR4D0BWP7T port map(A1 => VGA_l052_n_64, A2 => VGA_l052_n_57, A3 => VGA_l052_n_28, A4 => VGA_l052_n_29, ZN => VGA_l052_n_70);
  VGA_l052_g2494 : AOI211D0BWP7T port map(A1 => VGA_l052_n_7, A2 => VGA_l052_n_10, B => VGA_l052_n_66, C => VGA_l052_n_51, ZN => VGA_l052_n_69);
  VGA_l052_g2495 : NR4D0BWP7T port map(A1 => VGA_l052_n_61, A2 => VGA_l052_n_63, A3 => VGA_l052_n_53, A4 => VGA_l052_n_57, ZN => VGA_l052_n_68);
  VGA_l052_g2496 : OAI31D0BWP7T port map(A1 => VGA_l052_n_15, A2 => VGA_l052_n_34, A3 => VGA_l052_n_60, B => VGA_l052_n_65, ZN => VGA_l052_n_67);
  VGA_l052_g2497 : AOI22D0BWP7T port map(A1 => VGA_l052_n_62, A2 => VGA_l052_n_50, B1 => VGA_l052_n_33, B2 => VGA_l052_n_9, ZN => VGA_l052_n_66);
  VGA_l052_g2498 : OA32D0BWP7T port map(A1 => VGA_l052_n_20, A2 => VGA_l052_n_33, A3 => VGA_l052_n_1, B1 => VGA_l052_n_60, B2 => VGA_l052_n_58, Z => VGA_l052_n_65);
  VGA_l052_g2499 : OR3D0BWP7T port map(A1 => VGA_l052_n_30, A2 => VGA_l052_n_52, A3 => VGA_l052_n_63, Z => VGA_l052_n_64);
  VGA_l052_g2500 : OAI211D0BWP7T port map(A1 => VGA_l052_n_5, A2 => VGA_l052_n_11, B => VGA_l052_n_45, C => VGA_l052_n_19, ZN => VGA_l052_n_62);
  VGA_l052_g2501 : OAI221D0BWP7T port map(A1 => VGA_l052_n_35, A2 => VGA_l052_n_22, B1 => VGA_l052_n_16, B2 => VGA_l052_n_26, C => VGA_l052_n_48, ZN => VGA_l052_n_61);
  VGA_l052_g2502 : OAI211D0BWP7T port map(A1 => VGA_l052_n_18, A2 => VGA_l052_n_38, B => VGA_l052_n_46, C => VGA_l052_n_54, ZN => VGA_l052_n_63);
  VGA_l052_g2503 : MOAI22D0BWP7T port map(A1 => VGA_l052_n_25, A2 => y_pos_b2(1), B1 => VGA_l052_n_47, B2 => y_pos_b2(1), ZN => VGA_l052_n_59);
  VGA_l052_g2504 : OAI211D0BWP7T port map(A1 => VGA_l052_n_11, A2 => VGA_l052_n_36, B => VGA_l052_n_43, C => VGA_l052_n_44, ZN => VGA_l052_n_58);
  VGA_l052_g2505 : AO21D0BWP7T port map(A1 => VGA_l052_n_33, A2 => VGA_l052_n_20, B => VGA_l052_n_1, Z => VGA_l052_n_60);
  VGA_l052_g2506 : AOI22D0BWP7T port map(A1 => VGA_l052_n_30, A2 => VGA_l052_n_12, B1 => VGA_l052_n_41, B2 => VGA_y(1), ZN => VGA_l052_n_56);
  VGA_l052_g2507 : AOI22D0BWP7T port map(A1 => VGA_l052_n_37, A2 => VGA_l052_n_13, B1 => VGA_l052_n_2, B2 => x_pos_b2(8), ZN => VGA_l052_n_55);
  VGA_l052_g2508 : MAOI22D0BWP7T port map(A1 => VGA_l052_n_21, A2 => VGA_y(9), B1 => VGA_l052_n_21, B2 => VGA_y(9), ZN => VGA_l052_n_54);
  VGA_l052_g2509 : MOAI22D0BWP7T port map(A1 => VGA_l052_n_28, A2 => VGA_l052_n_14, B1 => VGA_l052_n_28, B2 => VGA_l052_n_14, ZN => VGA_l052_n_53);
  VGA_l052_g2510 : MAOI22D0BWP7T port map(A1 => VGA_l052_n_31, A2 => VGA_l052_n_23, B1 => VGA_l052_n_31, B2 => VGA_l052_n_23, ZN => VGA_l052_n_57);
  VGA_l052_g2511 : MOAI22D0BWP7T port map(A1 => VGA_l052_n_26, A2 => VGA_y(5), B1 => VGA_l052_n_26, B2 => VGA_y(5), ZN => VGA_l052_n_52);
  VGA_l052_g2512 : OAI22D0BWP7T port map(A1 => VGA_l052_n_40, A2 => VGA_l052_n_6, B1 => VGA_l052_n_32, B2 => VGA_l052_n_8, ZN => VGA_l052_n_51);
  VGA_l052_g2513 : MAOI22D0BWP7T port map(A1 => VGA_l052_n_34, A2 => VGA_l052_n_24, B1 => VGA_l052_n_33, B2 => VGA_l052_n_9, ZN => VGA_l052_n_50);
  VGA_l052_g2514 : MAOI22D0BWP7T port map(A1 => VGA_l052_n_32, A2 => VGA_l052_n_8, B1 => VGA_l052_n_7, B2 => VGA_l052_n_10, ZN => VGA_l052_n_49);
  VGA_l052_g2515 : AOI22D0BWP7T port map(A1 => VGA_l052_n_26, A2 => VGA_l052_n_16, B1 => VGA_l052_n_35, B2 => VGA_l052_n_22, ZN => VGA_l052_n_48);
  VGA_l052_g2517 : ND2D0BWP7T port map(A1 => VGA_l052_n_38, A2 => VGA_l052_n_18, ZN => VGA_l052_n_46);
  VGA_l052_g2518 : IND2D0BWP7T port map(A1 => VGA_l052_n_34, B1 => VGA_l052_n_15, ZN => VGA_l052_n_45);
  VGA_l052_g2519 : NR2D0BWP7T port map(A1 => VGA_l052_n_41, A2 => VGA_y(1), ZN => VGA_l052_n_47);
  VGA_l052_g2520 : ND2D0BWP7T port map(A1 => VGA_l052_n_34, A2 => VGA_l052_n_15, ZN => VGA_l052_n_44);
  VGA_l052_g2521 : AO21D0BWP7T port map(A1 => VGA_l052_n_36, A2 => VGA_l052_n_19, B => VGA_l052_n_5, Z => VGA_l052_n_43);
  VGA_l052_g2522 : CKXOR2D0BWP7T port map(A1 => VGA_y(0), A2 => VGA_l052_n_27, Z => VGA_l052_n_42);
  VGA_l052_g2525 : CKND1BWP7T port map(I => VGA_l052_n_25, ZN => VGA_l052_n_41);
  VGA_l052_g2526 : MOAI22D0BWP7T port map(A1 => VGA_x(6), A2 => x_pos_b2(6), B1 => VGA_x(6), B2 => x_pos_b2(6), ZN => VGA_l052_n_40);
  VGA_l052_g2527 : OA21D0BWP7T port map(A1 => VGA_l052_n_4, A2 => VGA_draw_count2(1), B => VGA_l052_n_17, Z => VGA_l052_n_39);
  VGA_l052_g2528 : MOAI22D0BWP7T port map(A1 => VGA_y(8), A2 => y_pos_b2(8), B1 => VGA_y(8), B2 => y_pos_b2(8), ZN => VGA_l052_n_38);
  VGA_l052_g2529 : MOAI22D0BWP7T port map(A1 => VGA_x(5), A2 => x_pos_b2(5), B1 => VGA_x(5), B2 => x_pos_b2(5), ZN => VGA_l052_n_37);
  VGA_l052_g2530 : AN2D1BWP7T port map(A1 => VGA_l052_n_15, A2 => VGA_l052_n_24, Z => VGA_l052_n_36);
  VGA_l052_g2531 : AO21D0BWP7T port map(A1 => VGA_l052_n_3, A2 => y_pos_b2(5), B => VGA_l052_n_16, Z => VGA_l052_n_35);
  VGA_l052_g2532 : MOAI22D0BWP7T port map(A1 => VGA_x(3), A2 => x_pos_b2(3), B1 => VGA_x(3), B2 => x_pos_b2(3), ZN => VGA_l052_n_34);
  VGA_l052_g2533 : MAOI22D0BWP7T port map(A1 => VGA_x(4), A2 => x_pos_b2(4), B1 => VGA_x(4), B2 => x_pos_b2(4), ZN => VGA_l052_n_33);
  VGA_l052_g2535 : MAOI22D0BWP7T port map(A1 => VGA_x(7), A2 => x_pos_b2(7), B1 => VGA_x(7), B2 => x_pos_b2(7), ZN => VGA_l052_n_32);
  VGA_l052_g2536 : MAOI22D0BWP7T port map(A1 => VGA_y(7), A2 => y_pos_b2(7), B1 => VGA_y(7), B2 => y_pos_b2(7), ZN => VGA_l052_n_31);
  VGA_l052_g2537 : MAOI22D0BWP7T port map(A1 => VGA_y(3), A2 => y_pos_b2(3), B1 => VGA_y(3), B2 => y_pos_b2(3), ZN => VGA_l052_n_30);
  VGA_l052_g2538 : MAOI22D0BWP7T port map(A1 => VGA_y(0), A2 => y_pos_b2(0), B1 => VGA_y(0), B2 => y_pos_b2(0), ZN => VGA_l052_n_29);
  VGA_l052_g2539 : MAOI22D0BWP7T port map(A1 => VGA_y(4), A2 => y_pos_b2(4), B1 => VGA_y(4), B2 => y_pos_b2(4), ZN => VGA_l052_n_28);
  VGA_l052_g2540 : MOAI22D0BWP7T port map(A1 => VGA_y(1), A2 => y_pos_b2(1), B1 => VGA_y(1), B2 => y_pos_b2(1), ZN => VGA_l052_n_27);
  VGA_l052_g2541 : MAOI22D0BWP7T port map(A1 => VGA_y(6), A2 => y_pos_b2(6), B1 => VGA_y(6), B2 => y_pos_b2(6), ZN => VGA_l052_n_26);
  VGA_l052_g2542 : MOAI22D0BWP7T port map(A1 => VGA_y(2), A2 => y_pos_b2(2), B1 => VGA_y(2), B2 => y_pos_b2(2), ZN => VGA_l052_n_25);
  VGA_l052_g2543 : IND2D0BWP7T port map(A1 => x_pos_b2(2), B1 => VGA_x(2), ZN => VGA_l052_n_24);
  VGA_l052_g2544 : INR2D0BWP7T port map(A1 => y_pos_b2(6), B1 => VGA_y(6), ZN => VGA_l052_n_23);
  VGA_l052_g2545 : INR2D0BWP7T port map(A1 => y_pos_b2(4), B1 => VGA_y(4), ZN => VGA_l052_n_22);
  VGA_l052_g2546 : IND2D0BWP7T port map(A1 => VGA_y(8), B1 => y_pos_b2(8), ZN => VGA_l052_n_21);
  VGA_l052_g2547 : INR2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_b2(3), ZN => VGA_l052_n_20);
  VGA_l052_g2548 : IND2D0BWP7T port map(A1 => x_pos_b2(1), B1 => VGA_x(1), ZN => VGA_l052_n_19);
  VGA_l052_g2549 : INR2D0BWP7T port map(A1 => y_pos_b2(7), B1 => VGA_y(7), ZN => VGA_l052_n_18);
  VGA_l052_g2550 : OR2D0BWP7T port map(A1 => VGA_draw_count2(2), A2 => VGA_draw_count2(1), Z => VGA_l052_n_17);
  VGA_l052_g2551 : NR2D0BWP7T port map(A1 => VGA_l052_n_3, A2 => y_pos_b2(5), ZN => VGA_l052_n_16);
  VGA_l052_g2552 : IND2D0BWP7T port map(A1 => VGA_x(2), B1 => x_pos_b2(2), ZN => VGA_l052_n_15);
  VGA_l052_g2553 : IND2D0BWP7T port map(A1 => VGA_y(3), B1 => y_pos_b2(3), ZN => VGA_l052_n_14);
  VGA_l052_g2554 : INR2D0BWP7T port map(A1 => x_pos_b2(4), B1 => VGA_x(4), ZN => VGA_l052_n_13);
  VGA_l052_g2555 : IND2D0BWP7T port map(A1 => VGA_y(2), B1 => y_pos_b2(2), ZN => VGA_l052_n_12);
  VGA_l052_g2556 : INR2D0BWP7T port map(A1 => x_pos_b2(1), B1 => VGA_x(1), ZN => VGA_l052_n_11);
  VGA_l052_g2557 : IND2D0BWP7T port map(A1 => x_pos_b2(8), B1 => VGA_x(8), ZN => VGA_l052_n_10);
  VGA_l052_g2558 : IND2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_b2(3), ZN => VGA_l052_n_9);
  VGA_l052_g2559 : INR2D0BWP7T port map(A1 => VGA_x(6), B1 => x_pos_b2(6), ZN => VGA_l052_n_8);
  VGA_l052_g2560 : INR2D0BWP7T port map(A1 => x_pos_b2(7), B1 => VGA_x(7), ZN => VGA_l052_n_7);
  VGA_l052_g2561 : IND2D0BWP7T port map(A1 => VGA_x(5), B1 => x_pos_b2(5), ZN => VGA_l052_n_6);
  VGA_l052_g2562 : IND2D0BWP7T port map(A1 => x_pos_b2(0), B1 => VGA_x(0), ZN => VGA_l052_n_5);
  VGA_l052_g2563 : CKND1BWP7T port map(I => VGA_draw_count2(0), ZN => VGA_l052_n_4);
  VGA_l052_g2564 : CKND1BWP7T port map(I => VGA_y(5), ZN => VGA_l052_n_3);
  VGA_l052_g2565 : CKND1BWP7T port map(I => VGA_x(8), ZN => VGA_l052_n_2);
  VGA_l052_g2 : MOAI22D0BWP7T port map(A1 => VGA_l052_n_37, A2 => VGA_l052_n_13, B1 => VGA_l052_n_40, B2 => VGA_l052_n_6, ZN => VGA_l052_n_1);
  VGA_l052_g2566 : INR4D0BWP7T port map(A1 => VGA_l052_n_29, B1 => VGA_l052_n_71, B2 => VGA_l052_n_59, B3 => VGA_l052_n_42, ZN => VGA_l052_n_0);
  VGA_l053_g2479 : AO31D0BWP7T port map(A1 => VGA_l053_n_77, A2 => VGA_l053_n_76, A3 => VGA_draw_count3(0), B => VGA_b3, Z => VGA_g3);
  VGA_l053_g2480 : OA21D0BWP7T port map(A1 => VGA_l053_n_79, A2 => VGA_l053_n_39, B => VGA_enable3, Z => VGA_r3);
  VGA_l053_g2481 : AO32D0BWP7T port map(A1 => VGA_l053_n_77, A2 => VGA_l053_n_76, A3 => VGA_l053_n_17, B1 => VGA_l053_n_78, B2 => VGA_l053_n_39, Z => VGA_b3);
  VGA_l053_g2482 : IND2D0BWP7T port map(A1 => VGA_l053_n_77, B1 => VGA_l053_n_75, ZN => VGA_enable3);
  VGA_l053_g2483 : MOAI22D0BWP7T port map(A1 => VGA_l053_n_4, A2 => VGA_draw_count3(2), B1 => VGA_l053_n_76, B2 => VGA_l053_n_73, ZN => VGA_l053_n_79);
  VGA_l053_g2484 : ND2D0BWP7T port map(A1 => VGA_l053_n_76, A2 => VGA_l053_n_75, ZN => VGA_l053_n_78);
  VGA_l053_g2485 : IAO21D0BWP7T port map(A1 => VGA_l053_n_74, A2 => VGA_l053_n_0, B => VGA_l053_n_72, ZN => VGA_l053_n_77);
  VGA_l053_g2486 : IND2D0BWP7T port map(A1 => VGA_l053_n_72, B1 => VGA_l053_n_74, ZN => VGA_l053_n_76);
  VGA_l053_g2487 : OR2D0BWP7T port map(A1 => VGA_l053_n_73, A2 => VGA_l053_n_72, Z => VGA_l053_n_75);
  VGA_l053_g2489 : NR4D0BWP7T port map(A1 => VGA_l053_n_71, A2 => VGA_l053_n_47, A3 => VGA_l053_n_29, A4 => VGA_l053_n_27, ZN => VGA_l053_n_74);
  VGA_l053_g2490 : ND4D0BWP7T port map(A1 => VGA_l053_n_70, A2 => VGA_l053_n_35, A3 => VGA_l053_n_27, A4 => VGA_l053_n_25, ZN => VGA_l053_n_73);
  VGA_l053_g2491 : ND4D0BWP7T port map(A1 => VGA_l053_n_67, A2 => VGA_l053_n_69, A3 => VGA_l053_n_55, A4 => VGA_l053_n_49, ZN => VGA_l053_n_72);
  VGA_l053_g2492 : OAI211D0BWP7T port map(A1 => VGA_l053_n_12, A2 => VGA_l053_n_30, B => VGA_l053_n_68, C => VGA_l053_n_56, ZN => VGA_l053_n_71);
  VGA_l053_g2493 : NR4D0BWP7T port map(A1 => VGA_l053_n_64, A2 => VGA_l053_n_57, A3 => VGA_l053_n_28, A4 => VGA_l053_n_29, ZN => VGA_l053_n_70);
  VGA_l053_g2494 : AOI211D0BWP7T port map(A1 => VGA_l053_n_7, A2 => VGA_l053_n_10, B => VGA_l053_n_66, C => VGA_l053_n_51, ZN => VGA_l053_n_69);
  VGA_l053_g2495 : NR4D0BWP7T port map(A1 => VGA_l053_n_61, A2 => VGA_l053_n_63, A3 => VGA_l053_n_53, A4 => VGA_l053_n_57, ZN => VGA_l053_n_68);
  VGA_l053_g2496 : OAI31D0BWP7T port map(A1 => VGA_l053_n_15, A2 => VGA_l053_n_34, A3 => VGA_l053_n_60, B => VGA_l053_n_65, ZN => VGA_l053_n_67);
  VGA_l053_g2497 : AOI22D0BWP7T port map(A1 => VGA_l053_n_62, A2 => VGA_l053_n_50, B1 => VGA_l053_n_33, B2 => VGA_l053_n_9, ZN => VGA_l053_n_66);
  VGA_l053_g2498 : OA32D0BWP7T port map(A1 => VGA_l053_n_20, A2 => VGA_l053_n_33, A3 => VGA_l053_n_1, B1 => VGA_l053_n_60, B2 => VGA_l053_n_58, Z => VGA_l053_n_65);
  VGA_l053_g2499 : OR3D0BWP7T port map(A1 => VGA_l053_n_30, A2 => VGA_l053_n_52, A3 => VGA_l053_n_63, Z => VGA_l053_n_64);
  VGA_l053_g2500 : OAI211D0BWP7T port map(A1 => VGA_l053_n_5, A2 => VGA_l053_n_11, B => VGA_l053_n_45, C => VGA_l053_n_19, ZN => VGA_l053_n_62);
  VGA_l053_g2501 : OAI221D0BWP7T port map(A1 => VGA_l053_n_35, A2 => VGA_l053_n_22, B1 => VGA_l053_n_16, B2 => VGA_l053_n_26, C => VGA_l053_n_48, ZN => VGA_l053_n_61);
  VGA_l053_g2502 : OAI211D0BWP7T port map(A1 => VGA_l053_n_18, A2 => VGA_l053_n_38, B => VGA_l053_n_46, C => VGA_l053_n_54, ZN => VGA_l053_n_63);
  VGA_l053_g2503 : MOAI22D0BWP7T port map(A1 => VGA_l053_n_25, A2 => y_pos_b3(1), B1 => VGA_l053_n_47, B2 => y_pos_b3(1), ZN => VGA_l053_n_59);
  VGA_l053_g2504 : OAI211D0BWP7T port map(A1 => VGA_l053_n_11, A2 => VGA_l053_n_36, B => VGA_l053_n_43, C => VGA_l053_n_44, ZN => VGA_l053_n_58);
  VGA_l053_g2505 : AO21D0BWP7T port map(A1 => VGA_l053_n_33, A2 => VGA_l053_n_20, B => VGA_l053_n_1, Z => VGA_l053_n_60);
  VGA_l053_g2506 : AOI22D0BWP7T port map(A1 => VGA_l053_n_30, A2 => VGA_l053_n_12, B1 => VGA_l053_n_41, B2 => VGA_y(1), ZN => VGA_l053_n_56);
  VGA_l053_g2507 : AOI22D0BWP7T port map(A1 => VGA_l053_n_37, A2 => VGA_l053_n_13, B1 => VGA_l053_n_2, B2 => x_pos_b3(8), ZN => VGA_l053_n_55);
  VGA_l053_g2508 : MAOI22D0BWP7T port map(A1 => VGA_l053_n_21, A2 => VGA_y(9), B1 => VGA_l053_n_21, B2 => VGA_y(9), ZN => VGA_l053_n_54);
  VGA_l053_g2509 : MOAI22D0BWP7T port map(A1 => VGA_l053_n_28, A2 => VGA_l053_n_14, B1 => VGA_l053_n_28, B2 => VGA_l053_n_14, ZN => VGA_l053_n_53);
  VGA_l053_g2510 : MAOI22D0BWP7T port map(A1 => VGA_l053_n_31, A2 => VGA_l053_n_23, B1 => VGA_l053_n_31, B2 => VGA_l053_n_23, ZN => VGA_l053_n_57);
  VGA_l053_g2511 : MOAI22D0BWP7T port map(A1 => VGA_l053_n_26, A2 => VGA_y(5), B1 => VGA_l053_n_26, B2 => VGA_y(5), ZN => VGA_l053_n_52);
  VGA_l053_g2512 : OAI22D0BWP7T port map(A1 => VGA_l053_n_40, A2 => VGA_l053_n_6, B1 => VGA_l053_n_32, B2 => VGA_l053_n_8, ZN => VGA_l053_n_51);
  VGA_l053_g2513 : MAOI22D0BWP7T port map(A1 => VGA_l053_n_34, A2 => VGA_l053_n_24, B1 => VGA_l053_n_33, B2 => VGA_l053_n_9, ZN => VGA_l053_n_50);
  VGA_l053_g2514 : MAOI22D0BWP7T port map(A1 => VGA_l053_n_32, A2 => VGA_l053_n_8, B1 => VGA_l053_n_7, B2 => VGA_l053_n_10, ZN => VGA_l053_n_49);
  VGA_l053_g2515 : AOI22D0BWP7T port map(A1 => VGA_l053_n_26, A2 => VGA_l053_n_16, B1 => VGA_l053_n_35, B2 => VGA_l053_n_22, ZN => VGA_l053_n_48);
  VGA_l053_g2517 : ND2D0BWP7T port map(A1 => VGA_l053_n_38, A2 => VGA_l053_n_18, ZN => VGA_l053_n_46);
  VGA_l053_g2518 : IND2D0BWP7T port map(A1 => VGA_l053_n_34, B1 => VGA_l053_n_15, ZN => VGA_l053_n_45);
  VGA_l053_g2519 : NR2D0BWP7T port map(A1 => VGA_l053_n_41, A2 => VGA_y(1), ZN => VGA_l053_n_47);
  VGA_l053_g2520 : ND2D0BWP7T port map(A1 => VGA_l053_n_34, A2 => VGA_l053_n_15, ZN => VGA_l053_n_44);
  VGA_l053_g2521 : AO21D0BWP7T port map(A1 => VGA_l053_n_36, A2 => VGA_l053_n_19, B => VGA_l053_n_5, Z => VGA_l053_n_43);
  VGA_l053_g2522 : CKXOR2D0BWP7T port map(A1 => VGA_y(0), A2 => VGA_l053_n_27, Z => VGA_l053_n_42);
  VGA_l053_g2525 : CKND1BWP7T port map(I => VGA_l053_n_25, ZN => VGA_l053_n_41);
  VGA_l053_g2526 : MOAI22D0BWP7T port map(A1 => VGA_x(6), A2 => x_pos_b3(6), B1 => VGA_x(6), B2 => x_pos_b3(6), ZN => VGA_l053_n_40);
  VGA_l053_g2527 : OA21D0BWP7T port map(A1 => VGA_l053_n_4, A2 => VGA_draw_count3(1), B => VGA_l053_n_17, Z => VGA_l053_n_39);
  VGA_l053_g2528 : MOAI22D0BWP7T port map(A1 => VGA_y(8), A2 => y_pos_b3(8), B1 => VGA_y(8), B2 => y_pos_b3(8), ZN => VGA_l053_n_38);
  VGA_l053_g2529 : MOAI22D0BWP7T port map(A1 => VGA_x(5), A2 => x_pos_b3(5), B1 => VGA_x(5), B2 => x_pos_b3(5), ZN => VGA_l053_n_37);
  VGA_l053_g2530 : AN2D1BWP7T port map(A1 => VGA_l053_n_15, A2 => VGA_l053_n_24, Z => VGA_l053_n_36);
  VGA_l053_g2531 : AO21D0BWP7T port map(A1 => VGA_l053_n_3, A2 => y_pos_b3(5), B => VGA_l053_n_16, Z => VGA_l053_n_35);
  VGA_l053_g2532 : MOAI22D0BWP7T port map(A1 => VGA_x(3), A2 => x_pos_b3(3), B1 => VGA_x(3), B2 => x_pos_b3(3), ZN => VGA_l053_n_34);
  VGA_l053_g2533 : MAOI22D0BWP7T port map(A1 => VGA_x(4), A2 => x_pos_b3(4), B1 => VGA_x(4), B2 => x_pos_b3(4), ZN => VGA_l053_n_33);
  VGA_l053_g2535 : MAOI22D0BWP7T port map(A1 => VGA_x(7), A2 => x_pos_b3(7), B1 => VGA_x(7), B2 => x_pos_b3(7), ZN => VGA_l053_n_32);
  VGA_l053_g2536 : MAOI22D0BWP7T port map(A1 => VGA_y(7), A2 => y_pos_b3(7), B1 => VGA_y(7), B2 => y_pos_b3(7), ZN => VGA_l053_n_31);
  VGA_l053_g2537 : MAOI22D0BWP7T port map(A1 => VGA_y(3), A2 => y_pos_b3(3), B1 => VGA_y(3), B2 => y_pos_b3(3), ZN => VGA_l053_n_30);
  VGA_l053_g2538 : MAOI22D0BWP7T port map(A1 => VGA_y(0), A2 => y_pos_b3(0), B1 => VGA_y(0), B2 => y_pos_b3(0), ZN => VGA_l053_n_29);
  VGA_l053_g2539 : MAOI22D0BWP7T port map(A1 => VGA_y(4), A2 => y_pos_b3(4), B1 => VGA_y(4), B2 => y_pos_b3(4), ZN => VGA_l053_n_28);
  VGA_l053_g2540 : MOAI22D0BWP7T port map(A1 => VGA_y(1), A2 => y_pos_b3(1), B1 => VGA_y(1), B2 => y_pos_b3(1), ZN => VGA_l053_n_27);
  VGA_l053_g2541 : MAOI22D0BWP7T port map(A1 => VGA_y(6), A2 => y_pos_b3(6), B1 => VGA_y(6), B2 => y_pos_b3(6), ZN => VGA_l053_n_26);
  VGA_l053_g2542 : MOAI22D0BWP7T port map(A1 => VGA_y(2), A2 => y_pos_b3(2), B1 => VGA_y(2), B2 => y_pos_b3(2), ZN => VGA_l053_n_25);
  VGA_l053_g2543 : IND2D0BWP7T port map(A1 => x_pos_b3(2), B1 => VGA_x(2), ZN => VGA_l053_n_24);
  VGA_l053_g2544 : INR2D0BWP7T port map(A1 => y_pos_b3(6), B1 => VGA_y(6), ZN => VGA_l053_n_23);
  VGA_l053_g2545 : INR2D0BWP7T port map(A1 => y_pos_b3(4), B1 => VGA_y(4), ZN => VGA_l053_n_22);
  VGA_l053_g2546 : IND2D0BWP7T port map(A1 => VGA_y(8), B1 => y_pos_b3(8), ZN => VGA_l053_n_21);
  VGA_l053_g2547 : INR2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_b3(3), ZN => VGA_l053_n_20);
  VGA_l053_g2548 : IND2D0BWP7T port map(A1 => x_pos_b3(1), B1 => VGA_x(1), ZN => VGA_l053_n_19);
  VGA_l053_g2549 : INR2D0BWP7T port map(A1 => y_pos_b3(7), B1 => VGA_y(7), ZN => VGA_l053_n_18);
  VGA_l053_g2550 : OR2D0BWP7T port map(A1 => VGA_draw_count3(2), A2 => VGA_draw_count3(1), Z => VGA_l053_n_17);
  VGA_l053_g2551 : NR2D0BWP7T port map(A1 => VGA_l053_n_3, A2 => y_pos_b3(5), ZN => VGA_l053_n_16);
  VGA_l053_g2552 : IND2D0BWP7T port map(A1 => VGA_x(2), B1 => x_pos_b3(2), ZN => VGA_l053_n_15);
  VGA_l053_g2553 : IND2D0BWP7T port map(A1 => VGA_y(3), B1 => y_pos_b3(3), ZN => VGA_l053_n_14);
  VGA_l053_g2554 : INR2D0BWP7T port map(A1 => x_pos_b3(4), B1 => VGA_x(4), ZN => VGA_l053_n_13);
  VGA_l053_g2555 : IND2D0BWP7T port map(A1 => VGA_y(2), B1 => y_pos_b3(2), ZN => VGA_l053_n_12);
  VGA_l053_g2556 : INR2D0BWP7T port map(A1 => x_pos_b3(1), B1 => VGA_x(1), ZN => VGA_l053_n_11);
  VGA_l053_g2557 : IND2D0BWP7T port map(A1 => x_pos_b3(8), B1 => VGA_x(8), ZN => VGA_l053_n_10);
  VGA_l053_g2558 : IND2D0BWP7T port map(A1 => VGA_x(3), B1 => x_pos_b3(3), ZN => VGA_l053_n_9);
  VGA_l053_g2559 : INR2D0BWP7T port map(A1 => VGA_x(6), B1 => x_pos_b3(6), ZN => VGA_l053_n_8);
  VGA_l053_g2560 : INR2D0BWP7T port map(A1 => x_pos_b3(7), B1 => VGA_x(7), ZN => VGA_l053_n_7);
  VGA_l053_g2561 : IND2D0BWP7T port map(A1 => VGA_x(5), B1 => x_pos_b3(5), ZN => VGA_l053_n_6);
  VGA_l053_g2562 : IND2D0BWP7T port map(A1 => x_pos_b3(0), B1 => VGA_x(0), ZN => VGA_l053_n_5);
  VGA_l053_g2563 : CKND1BWP7T port map(I => VGA_draw_count3(0), ZN => VGA_l053_n_4);
  VGA_l053_g2564 : CKND1BWP7T port map(I => VGA_y(5), ZN => VGA_l053_n_3);
  VGA_l053_g2565 : CKND1BWP7T port map(I => VGA_x(8), ZN => VGA_l053_n_2);
  VGA_l053_g2 : MOAI22D0BWP7T port map(A1 => VGA_l053_n_37, A2 => VGA_l053_n_13, B1 => VGA_l053_n_40, B2 => VGA_l053_n_6, ZN => VGA_l053_n_1);
  VGA_l053_g2566 : INR4D0BWP7T port map(A1 => VGA_l053_n_29, B1 => VGA_l053_n_71, B2 => VGA_l053_n_59, B3 => VGA_l053_n_42, ZN => VGA_l053_n_0);
  Enemy_spawning_en61_decider_reg : DFQD1BWP7T port map(CP => clk, D => Enemy_spawning_en61_n_3, Q => spawn_or_not_e6);
  Enemy_spawning_en61_g143 : NR4D0BWP7T port map(A1 => Enemy_spawning_en61_n_2, A2 => Enemy_spawning_en61_n_1, A3 => Enemy_spawning_en61_n_0, A4 => e_6, ZN => Enemy_spawning_en61_n_3);
  Enemy_spawning_en61_g144 : ND4D0BWP7T port map(A1 => y_e_spawn_3(1), A2 => y_e_spawn_3(7), A3 => y_e_spawn_1(2), A4 => y_e_spawn_1(3), ZN => Enemy_spawning_en61_n_2);
  Enemy_spawning_en61_g145 : ND2D0BWP7T port map(A1 => y_e_spawn_4(7), A2 => y_e_spawn_2(3), ZN => Enemy_spawning_en61_n_1);
  Enemy_spawning_en61_g146 : ND2D0BWP7T port map(A1 => y_e_spawn_5(8), A2 => n_5, ZN => Enemy_spawning_en61_n_0);
  Collision_L1_range_state_out_reg_1 : DFQD1BWP7T port map(CP => clk, D => Collision_L1_n_479, Q => Collision_L1_range_state_out(1));
  Collision_L1_g3368 : AOI221D0BWP7T port map(A1 => Collision_L1_n_482, A2 => Collision_L1_n_4, B1 => Collision_L1_n_481, B2 => Collision_L1_n_484, C => reset, ZN => Collision_L1_n_479);
  Collision_L1_g3369 : INVD1BWP7T port map(I => Collision_L1_n_4, ZN => Collision_L1_n_483);
  Collision_L1_g3370 : INR4D0BWP7T port map(A1 => Collision_count_2_s(2), B1 => Collision_count_2_s(3), B2 => Collision_count_2_s(1), B3 => Collision_count_2_s(0), ZN => Collision_L1_n_4);
  Collision_L1_g3371 : OA31D0BWP7T port map(A1 => Collision_count_2_s(1), A2 => Collision_count_2_s(2), A3 => Collision_count_2_s(0), B => Collision_count_2_s(3), Z => Collision_L1_n_481);
  Collision_L1_g3373 : OAI22D0BWP7T port map(A1 => Collision_L1_n_500, A2 => Collision_count_1_s(1), B1 => Collision_count_1_s(3), B2 => Collision_count_1_s(2), ZN => Collision_start_value_s(0));
  Collision_L1_g3374 : OA21D0BWP7T port map(A1 => Collision_L1_n_501, A2 => Collision_count_1_s(0), B => Collision_count_1_s(3), Z => Collision_L1_n_482);
  Collision_L1_g3376 : NR2D0BWP7T port map(A1 => Collision_L1_n_500, A2 => Collision_L1_n_502, ZN => Collision_L1_n_484);
  Collision_L1_g3377 : IND2D0BWP7T port map(A1 => Collision_enable_s, B1 => Collision_L1_state(0), ZN => Collision_reset_2_s);
  Collision_L1_g3378 : NR2D0BWP7T port map(A1 => Collision_count_1_s(3), A2 => Collision_count_1_s(2), ZN => Collision_start_value_s(3));
  Collision_L1_g3379 : IND2D0BWP7T port map(A1 => Collision_count_1_s(0), B1 => Collision_L1_n_476, ZN => Collision_L1_n_500);
  Collision_L1_g3380 : IND2D0BWP7T port map(A1 => Collision_count_1_s(1), B1 => Collision_count_1_s(2), ZN => Collision_L1_n_502);
  Collision_L1_g3381 : IND2D0BWP7T port map(A1 => Collision_count_1_s(0), B1 => Collision_count_1_s(3), ZN => Collision_L1_n_503);
  Collision_L1_g3382 : OR2D0BWP7T port map(A1 => Collision_count_1_s(2), A2 => Collision_count_1_s(1), Z => Collision_L1_n_501);
  Collision_L1_g3383 : INVD0BWP7T port map(I => Collision_count_1_s(3), ZN => Collision_L1_n_476);
  Collision_L1_col_reg_0 : DFQD1BWP7T port map(CP => clk, D => Collision_L1_n_238, Q => collision_output_vector(0));
  Collision_L1_col_reg_1 : DFQD1BWP7T port map(CP => clk, D => Collision_L1_n_245, Q => collision_output_vector(1));
  Collision_L1_col_reg_2 : DFQD1BWP7T port map(CP => clk, D => Collision_L1_n_240, Q => collision_output_vector(2));
  Collision_L1_col_reg_4 : DFQD1BWP7T port map(CP => clk, D => Collision_L1_n_246, Q => collision_output_vector(4));
  Collision_L1_col_reg_9 : DFQD1BWP7T port map(CP => clk, D => Collision_L1_n_239, Q => collision_output_vector(9));
  Collision_L1_col_reg_10 : DFQD1BWP7T port map(CP => clk, D => Collision_L1_n_244, Q => collision_output_vector(10));
  Collision_L1_col_reg_11 : DFQD1BWP7T port map(CP => clk, D => Collision_L1_n_243, Q => collision_output_vector(11));
  Collision_L1_col_reg_12 : DFQD1BWP7T port map(CP => clk, D => Collision_L1_n_242, Q => collision_output_vector(12));
  Collision_L1_col_reg_13 : DFQD1BWP7T port map(CP => clk, D => Collision_L1_n_241, Q => collision_output_vector(13));
  Collision_L1_col_reg_14 : DFQD1BWP7T port map(CP => clk, D => Collision_L1_n_250, Q => collision_output_vector(14));
  Collision_L1_state_reg_0 : DFND1BWP7T port map(CPN => clk, D => Collision_L1_n_475, Q => Collision_L1_state(0), QN => Collision_L1_n_2);
  Collision_L1_state_reg_1 : DFND1BWP7T port map(CPN => clk, D => Collision_L1_n_474, Q => Collision_enable_s, QN => UNCONNECTED1);
  Collision_L1_state_reg_2 : DFND1BWP7T port map(CPN => clk, D => Collision_L1_n_216, Q => Collision_L1_state(2), QN => UNCONNECTED2);
  Collision_L1_g14031 : OAI222D0BWP7T port map(A1 => Collision_L1_n_473, A2 => Collision_L1_n_54, B1 => Collision_L1_n_21, B2 => Collision_L1_n_35, C1 => Collision_L1_n_50, C2 => Collision_L1_n_16, ZN => Collision_L1_n_475);
  Collision_L1_g14032 : IAO21D0BWP7T port map(A1 => Collision_L1_n_473, A2 => Collision_L1_n_168, B => Collision_L1_n_54, ZN => Collision_L1_n_474);
  Collision_L1_g14033 : ND2D0BWP7T port map(A1 => Collision_L1_n_472, A2 => Collision_L1_n_438, ZN => Collision_L1_n_473);
  Collision_L1_g14034 : AOI221D0BWP7T port map(A1 => Collision_L1_n_382, A2 => Collision_L1_n_269, B1 => Collision_L1_n_389, B2 => Collision_L1_n_291, C => Collision_L1_n_471, ZN => Collision_L1_n_472);
  Collision_L1_g14035 : INR4D0BWP7T port map(A1 => Collision_L1_n_455, B1 => Collision_L1_n_467, B2 => Collision_L1_n_464, B3 => Collision_L1_n_470, ZN => Collision_L1_n_471);
  Collision_L1_g14036 : OAI21D0BWP7T port map(A1 => Collision_L1_n_436, A2 => Collision_L1_n_297, B => Collision_L1_n_469, ZN => Collision_L1_n_470);
  Collision_L1_g14037 : AO221D0BWP7T port map(A1 => Collision_L1_n_459, A2 => Collision_L1_n_298, B1 => Collision_L1_n_465, B2 => Collision_L1_n_433, C => Collision_L1_n_468, Z => Collision_L1_n_469);
  Collision_L1_g14038 : OAI221D0BWP7T port map(A1 => Collision_L1_n_462, A2 => Collision_L1_n_411, B1 => Collision_L1_n_296, B2 => Collision_L1_n_451, C => Collision_L1_n_466, ZN => Collision_L1_n_468);
  Collision_L1_g14039 : AOI221D0BWP7T port map(A1 => Collision_L1_n_456, A2 => Collision_L1_n_432, B1 => Collision_L1_n_436, B2 => Collision_L1_n_297, C => Collision_L1_n_463, ZN => Collision_L1_n_467);
  Collision_L1_g14040 : AOI33D0BWP7T port map(A1 => Collision_L1_n_461, A2 => Collision_L1_n_428, A3 => Collision_L1_n_303, B1 => Collision_L1_n_457, B2 => Collision_L1_n_443, B3 => Collision_L1_n_301, ZN => Collision_L1_n_466);
  Collision_L1_g14041 : OAI31D0BWP7T port map(A1 => Collision_L1_n_411, A2 => Collision_L1_n_441, A3 => Collision_L1_n_460, B => Collision_L1_n_462, ZN => Collision_L1_n_465);
  Collision_L1_g14042 : OAI211D0BWP7T port map(A1 => Collision_L1_n_298, A2 => Collision_L1_n_459, B => Collision_L1_n_450, C => Collision_L1_n_60, ZN => Collision_L1_n_464);
  Collision_L1_g14043 : OAI221D0BWP7T port map(A1 => Collision_L1_n_454, A2 => Collision_L1_n_396, B1 => Collision_L1_n_312, B2 => Collision_L1_n_446, C => Collision_L1_n_458, ZN => Collision_L1_n_463);
  Collision_L1_g14044 : IND3D0BWP7T port map(A1 => Collision_L1_n_441, B1 => Collision_L1_n_305, B2 => Collision_L1_n_461, ZN => Collision_L1_n_462);
  Collision_L1_g14045 : CKND1BWP7T port map(I => Collision_L1_n_460, ZN => Collision_L1_n_461);
  Collision_L1_g14046 : OAI21D0BWP7T port map(A1 => Collision_L1_n_443, A2 => Collision_L1_n_301, B => Collision_L1_n_457, ZN => Collision_L1_n_460);
  Collision_L1_g14047 : AOI33D0BWP7T port map(A1 => Collision_L1_n_453, A2 => Collision_L1_n_416, A3 => Collision_L1_n_295, B1 => Collision_L1_n_449, B2 => Collision_L1_n_442, B3 => Collision_L1_n_310, ZN => Collision_L1_n_458);
  Collision_L1_g14048 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_448, A2 => Collision_L1_n_278, B1 => Collision_L1_n_448, B2 => Collision_L1_n_278, ZN => Collision_L1_n_459);
  Collision_L1_g14049 : ND2D0BWP7T port map(A1 => Collision_L1_n_451, A2 => Collision_L1_n_296, ZN => Collision_L1_n_457);
  Collision_L1_g14050 : OAI31D0BWP7T port map(A1 => Collision_L1_n_396, A2 => Collision_L1_n_427, A3 => Collision_L1_n_452, B => Collision_L1_n_454, ZN => Collision_L1_n_456);
  Collision_L1_g14051 : MAOI222D0BWP7T port map(A => Collision_L1_n_505, B => Collision_L1_n_297, C => Collision_L1_n_447, ZN => Collision_L1_n_455);
  Collision_L1_g14052 : IND3D0BWP7T port map(A1 => Collision_L1_n_427, B1 => Collision_L1_n_313, B2 => Collision_L1_n_453, ZN => Collision_L1_n_454);
  Collision_L1_g14053 : CKND1BWP7T port map(I => Collision_L1_n_452, ZN => Collision_L1_n_453);
  Collision_L1_g14054 : OAI21D0BWP7T port map(A1 => Collision_L1_n_442, A2 => Collision_L1_n_310, B => Collision_L1_n_449, ZN => Collision_L1_n_452);
  Collision_L1_g14055 : MAOI222D0BWP7T port map(A => Collision_L1_n_415, B => Collision_L1_n_298, C => Collision_L1_n_445, ZN => Collision_L1_n_450);
  Collision_L1_g14056 : OAI21D0BWP7T port map(A1 => Collision_L1_n_440, A2 => Collision_L1_n_291, B => Collision_L1_n_448, ZN => Collision_L1_n_451);
  Collision_L1_g14057 : ND2D0BWP7T port map(A1 => Collision_L1_n_446, A2 => Collision_L1_n_312, ZN => Collision_L1_n_449);
  Collision_L1_g14058 : ND2D0BWP7T port map(A1 => Collision_L1_n_440, A2 => Collision_L1_n_291, ZN => Collision_L1_n_448);
  Collision_L1_g14059 : AOI31D0BWP7T port map(A1 => Collision_L1_n_426, A2 => Collision_L1_n_431, A3 => Collision_L1_n_402, B => Collision_L1_n_444, ZN => Collision_L1_n_447);
  Collision_L1_g14060 : AOI221D0BWP7T port map(A1 => Collision_L1_n_429, A2 => Collision_L1_n_409, B1 => Collision_L1_n_429, B2 => Collision_L1_n_406, C => Collision_L1_n_437, ZN => Collision_L1_n_445);
  Collision_L1_g14061 : OAI21D0BWP7T port map(A1 => Collision_L1_n_439, A2 => Collision_L1_n_272, B => Collision_L1_n_425, ZN => Collision_L1_n_446);
  Collision_L1_g14062 : OAI31D0BWP7T port map(A1 => Collision_L1_n_310, A2 => Collision_L1_n_399, A3 => Collision_L1_n_420, B => Collision_L1_n_434, ZN => Collision_L1_n_444);
  Collision_L1_g14063 : AOI21D0BWP7T port map(A1 => Collision_L1_n_430, A2 => Collision_L1_n_290, B => Collision_L1_n_440, ZN => Collision_L1_n_443);
  Collision_L1_g14064 : HA1D0BWP7T port map(A => Collision_L1_n_265, B => Collision_L1_n_413, CO => Collision_L1_n_439, S => Collision_L1_n_442);
  Collision_L1_g14065 : AOI31D0BWP7T port map(A1 => Collision_L1_n_419, A2 => Collision_L1_n_506, A3 => Collision_L1_n_418, B => Collision_L1_n_393, ZN => Collision_L1_n_438);
  Collision_L1_g14066 : NR2D0BWP7T port map(A1 => Collision_L1_n_428, A2 => Collision_L1_n_303, ZN => Collision_L1_n_441);
  Collision_L1_g14067 : NR2D0BWP7T port map(A1 => Collision_L1_n_430, A2 => Collision_L1_n_290, ZN => Collision_L1_n_440);
  Collision_L1_g14068 : CKND1BWP7T port map(I => Collision_L1_n_435, ZN => Collision_L1_n_437);
  Collision_L1_g14069 : MAOI222D0BWP7T port map(A => Collision_L1_n_417, B => Collision_L1_n_296, C => Collision_L1_n_419, ZN => Collision_L1_n_435);
  Collision_L1_g14070 : AOI22D0BWP7T port map(A1 => Collision_L1_n_426, A2 => Collision_L1_n_424, B1 => Collision_L1_n_407, B2 => Collision_L1_n_312, ZN => Collision_L1_n_434);
  Collision_L1_g14071 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_425, A2 => Collision_L1_n_269, B1 => Collision_L1_n_425, B2 => Collision_L1_n_269, ZN => Collision_L1_n_436);
  Collision_L1_g14072 : MAOI222D0BWP7T port map(A => Collision_L1_n_371, B => Collision_L1_n_300, C => Collision_L1_n_404, ZN => Collision_L1_n_433);
  Collision_L1_g14073 : MAOI222D0BWP7T port map(A => Collision_L1_n_352, B => Collision_L1_n_311, C => Collision_L1_n_403, ZN => Collision_L1_n_432);
  Collision_L1_g14074 : AOI21D0BWP7T port map(A1 => Collision_L1_n_377, A2 => Collision_L1_n_313, B => Collision_L1_n_422, ZN => Collision_L1_n_431);
  Collision_L1_g14075 : OAI21D0BWP7T port map(A1 => Collision_L1_n_421, A2 => Collision_L1_range_state_out(0), B => Collision_L1_n_287, ZN => Collision_L1_n_430);
  Collision_L1_g14076 : OA21D0BWP7T port map(A1 => Collision_L1_n_419, A2 => Collision_L1_n_296, B => Collision_L1_n_423, Z => Collision_L1_n_429);
  Collision_L1_g14077 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_401, A2 => Collision_L1_n_325, B1 => Collision_L1_n_401, B2 => Collision_L1_n_325, ZN => Collision_L1_n_428);
  Collision_L1_g14078 : NR2D0BWP7T port map(A1 => Collision_L1_n_416, A2 => Collision_L1_n_295, ZN => Collision_L1_n_427);
  Collision_L1_g14079 : AOI21D0BWP7T port map(A1 => Collision_L1_n_399, A2 => Collision_L1_n_310, B => Collision_L1_n_420, ZN => Collision_L1_n_426);
  Collision_L1_g14080 : ND2D0BWP7T port map(A1 => Collision_L1_n_413, A2 => Collision_L1_n_316, ZN => Collision_L1_n_425);
  Collision_L1_g14081 : OAI22D0BWP7T port map(A1 => Collision_L1_n_408, A2 => Collision_L1_n_313, B1 => Collision_L1_n_390, B2 => Collision_L1_n_295, ZN => Collision_L1_n_424);
  Collision_L1_g14082 : AOI22D0BWP7T port map(A1 => Collision_L1_n_410, A2 => Collision_L1_n_301, B1 => Collision_L1_n_395, B2 => Collision_L1_n_303, ZN => Collision_L1_n_423);
  Collision_L1_g14083 : MAOI222D0BWP7T port map(A => Collision_L1_n_358, B => Collision_L1_n_311, C => Collision_L1_n_405, ZN => Collision_L1_n_422);
  Collision_L1_g14084 : CKND1BWP7T port map(I => Collision_L1_n_401, ZN => Collision_L1_n_421);
  Collision_L1_g14085 : OAI31D0BWP7T port map(A1 => Collision_L1_n_394, A2 => Collision_L1_n_376, A3 => Collision_L1_n_395, B => Collision_L1_n_410, ZN => Collision_L1_n_418);
  Collision_L1_g14086 : NR2D0BWP7T port map(A1 => Collision_L1_n_407, A2 => Collision_L1_n_312, ZN => Collision_L1_n_420);
  Collision_L1_g14087 : NR2D0BWP7T port map(A1 => Collision_L1_n_410, A2 => Collision_L1_n_301, ZN => Collision_L1_n_417);
  Collision_L1_g14088 : OAI221D0BWP7T port map(A1 => Collision_L1_n_392, A2 => Collision_L1_n_292, B1 => Collision_L1_n_291, B2 => Collision_L1_n_385, C => Collision_L1_n_12, ZN => Collision_L1_n_419);
  Collision_L1_g14089 : CKND1BWP7T port map(I => Collision_L1_n_506, ZN => Collision_L1_n_415);
  Collision_L1_g14091 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_383, A2 => Collision_L1_n_322, B1 => Collision_L1_n_383, B2 => Collision_L1_n_322, ZN => Collision_L1_n_416);
  Collision_L1_g14093 : AOI21D0BWP7T port map(A1 => Collision_L1_n_383, A2 => Collision_L1_n_3, B => Collision_L1_n_264, ZN => Collision_L1_n_413);
  Collision_L1_g14094 : AOI211D0BWP7T port map(A1 => Collision_L1_n_376, A2 => Collision_L1_n_305, B => Collision_L1_n_400, C => Collision_L1_n_381, ZN => Collision_L1_n_409);
  Collision_L1_g14095 : IND2D0BWP7T port map(A1 => Collision_L1_n_377, B1 => Collision_L1_n_402, ZN => Collision_L1_n_408);
  Collision_L1_g14096 : OAI21D0BWP7T port map(A1 => Collision_L1_n_368, A2 => Collision_L1_n_275, B => Collision_L1_n_401, ZN => Collision_L1_n_411);
  Collision_L1_g14097 : OA221D0BWP7T port map(A1 => Collision_L1_n_372, A2 => Collision_L1_n_290, B1 => Collision_L1_n_289, B2 => Collision_L1_n_375, C => Collision_L1_n_12, Z => Collision_L1_n_410);
  Collision_L1_g14098 : OAI22D0BWP7T port map(A1 => Collision_L1_n_395, A2 => Collision_L1_n_303, B1 => Collision_L1_n_376, B2 => Collision_L1_n_305, ZN => Collision_L1_n_406);
  Collision_L1_g14099 : MAOI222D0BWP7T port map(A => Collision_L1_n_349, B => Collision_L1_n_304, C => Collision_L1_n_370, ZN => Collision_L1_n_405);
  Collision_L1_g14100 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_363, A2 => Collision_L1_n_281, B1 => Collision_L1_n_387, B2 => Collision_L1_n_378, ZN => Collision_L1_n_404);
  Collision_L1_g14101 : OAI22D0BWP7T port map(A1 => Collision_L1_n_391, A2 => Collision_L1_n_273, B1 => Collision_L1_n_388, B2 => Collision_L1_n_272, ZN => Collision_L1_n_407);
  Collision_L1_g14102 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_362, A2 => Collision_L1_n_304, B1 => Collision_L1_n_386, B2 => Collision_L1_n_380, ZN => Collision_L1_n_403);
  Collision_L1_g14103 : AOI222D0BWP7T port map(A1 => Collision_L1_n_367, A2 => Collision_L1_n_300, B1 => Collision_L1_n_350, B2 => Collision_L1_n_282, C1 => Collision_L1_n_365, C2 => Collision_L1_n_359, ZN => Collision_L1_n_400);
  Collision_L1_g14104 : ND2D0BWP7T port map(A1 => Collision_L1_n_390, A2 => Collision_L1_n_295, ZN => Collision_L1_n_402);
  Collision_L1_g14105 : ND2D0BWP7T port map(A1 => Collision_L1_n_368, A2 => Collision_L1_n_275, ZN => Collision_L1_n_401);
  Collision_L1_g14108 : AOI22D0BWP7T port map(A1 => Collision_L1_n_374, A2 => Collision_L1_n_265, B1 => Collision_L1_n_373, B2 => Collision_L1_n_266, ZN => Collision_L1_n_399);
  Collision_L1_g14109 : AOI31D0BWP7T port map(A1 => Collision_L1_n_350, A2 => Collision_L1_n_323, A3 => Collision_L1_n_284, B => Collision_L1_n_367, ZN => Collision_L1_n_394);
  Collision_L1_g14110 : NR4D0BWP7T port map(A1 => Collision_L1_n_345, A2 => Collision_L1_n_264, A3 => Collision_L1_n_268, A4 => Collision_L1_n_294, ZN => Collision_L1_n_393);
  Collision_L1_g14111 : IAO21D0BWP7T port map(A1 => Collision_L1_n_369, A2 => Collision_L1_n_14, B => Collision_L1_n_332, ZN => Collision_L1_n_392);
  Collision_L1_g14112 : AOI21D0BWP7T port map(A1 => Collision_L1_n_366, A2 => Collision_L1_n_58, B => Collision_L1_n_334, ZN => Collision_L1_n_391);
  Collision_L1_g14113 : OAI21D0BWP7T port map(A1 => Collision_L1_n_342, A2 => Collision_L1_n_267, B => Collision_L1_n_383, ZN => Collision_L1_n_396);
  Collision_L1_g14114 : AOI32D0BWP7T port map(A1 => Collision_L1_n_343, A2 => Collision_L1_n_288, A3 => Collision_L1_n_58, B1 => Collision_L1_n_364, B2 => Collision_L1_n_287, ZN => Collision_L1_n_395);
  Collision_L1_g14115 : AOI211D0BWP7T port map(A1 => Collision_L1_n_351, A2 => Collision_L1_n_288, B => Collision_L1_n_290, C => Collision_L1_n_278, ZN => Collision_L1_n_389);
  Collision_L1_g14116 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_318, A2 => Collision_L1_n_34, B1 => Collision_L1_n_366, B2 => Collision_L1_n_14, ZN => Collision_L1_n_388);
  Collision_L1_g14117 : OAI22D0BWP7T port map(A1 => Collision_L1_n_363, A2 => Collision_L1_n_281, B1 => Collision_L1_n_328, B2 => Collision_L1_n_299, ZN => Collision_L1_n_387);
  Collision_L1_g14118 : OAI22D0BWP7T port map(A1 => Collision_L1_n_362, A2 => Collision_L1_n_304, B1 => Collision_L1_n_327, B2 => Collision_L1_n_302, ZN => Collision_L1_n_386);
  Collision_L1_g14119 : AOI22D0BWP7T port map(A1 => Collision_L1_n_369, A2 => Collision_L1_n_58, B1 => Collision_L1_n_319, B2 => Collision_L1_n_34, ZN => Collision_L1_n_385);
  Collision_L1_g14120 : AOI32D0BWP7T port map(A1 => Collision_L1_n_340, A2 => Collision_L1_n_264, A3 => Collision_L1_n_58, B1 => Collision_L1_n_361, B2 => Collision_L1_n_263, ZN => Collision_L1_n_390);
  Collision_L1_g14121 : OAI31D0BWP7T port map(A1 => Collision_L1_n_263, A2 => Collision_L1_n_267, A3 => Collision_L1_n_339, B => Collision_L1_n_316, ZN => Collision_L1_n_382);
  Collision_L1_g14122 : NR2D0BWP7T port map(A1 => Collision_L1_n_367, A2 => Collision_L1_n_300, ZN => Collision_L1_n_381);
  Collision_L1_g14123 : AOI211D0BWP7T port map(A1 => Collision_L1_n_327, A2 => Collision_L1_n_302, B => Collision_L1_n_307, C => Collision_L1_n_283, ZN => Collision_L1_n_380);
  Collision_L1_g14125 : AOI211D0BWP7T port map(A1 => Collision_L1_n_328, A2 => Collision_L1_n_299, B => Collision_L1_n_306, C => Collision_L1_n_285, ZN => Collision_L1_n_378);
  Collision_L1_g14127 : ND2D0BWP7T port map(A1 => Collision_L1_n_342, A2 => Collision_L1_n_267, ZN => Collision_L1_n_383);
  Collision_L1_g14128 : AOI22D0BWP7T port map(A1 => Collision_L1_n_353, A2 => Collision_L1_n_58, B1 => Collision_L1_n_287, B2 => Collision_L1_n_34, ZN => Collision_L1_n_375);
  Collision_L1_g14129 : OAI22D0BWP7T port map(A1 => Collision_L1_n_356, A2 => Collision_L1_n_14, B1 => Collision_L1_n_263, B2 => Collision_L1_n_59, ZN => Collision_L1_n_374);
  Collision_L1_g14130 : OAI22D0BWP7T port map(A1 => Collision_L1_n_355, A2 => Collision_L1_n_14, B1 => Collision_L1_n_264, B2 => Collision_L1_n_59, ZN => Collision_L1_n_373);
  Collision_L1_g14131 : AOI22D0BWP7T port map(A1 => Collision_L1_n_354, A2 => Collision_L1_n_58, B1 => Collision_L1_n_288, B2 => Collision_L1_n_34, ZN => Collision_L1_n_372);
  Collision_L1_g14132 : AO21D0BWP7T port map(A1 => Collision_L1_n_357, A2 => Collision_L1_n_274, B => Collision_L1_n_368, Z => Collision_L1_n_371);
  Collision_L1_g14133 : AOI32D0BWP7T port map(A1 => Collision_L1_n_321, A2 => Collision_L1_n_267, A3 => Collision_L1_n_58, B1 => Collision_L1_n_347, B2 => Collision_L1_n_268, ZN => Collision_L1_n_377);
  Collision_L1_g14134 : IOA21D0BWP7T port map(A1 => Collision_L1_n_337, A2 => Collision_L1_n_302, B => Collision_L1_n_360, ZN => Collision_L1_n_370);
  Collision_L1_g14135 : AOI32D0BWP7T port map(A1 => Collision_L1_n_331, A2 => Collision_L1_n_275, A3 => Collision_L1_n_58, B1 => Collision_L1_n_346, B2 => Collision_L1_n_276, ZN => Collision_L1_n_376);
  Collision_L1_g14136 : IND2D0BWP7T port map(A1 => Collision_L1_n_350, B1 => Collision_L1_n_281, ZN => Collision_L1_n_365);
  Collision_L1_g14137 : OAI21D0BWP7T port map(A1 => Collision_L1_n_343, A2 => Collision_L1_n_14, B => Collision_L1_n_59, ZN => Collision_L1_n_364);
  Collision_L1_g14138 : ND2D0BWP7T port map(A1 => Collision_L1_n_354, A2 => Collision_L1_n_290, ZN => Collision_L1_n_369);
  Collision_L1_g14139 : NR2D0BWP7T port map(A1 => Collision_L1_n_357, A2 => Collision_L1_n_274, ZN => Collision_L1_n_368);
  Collision_L1_g14140 : OAI31D0BWP7T port map(A1 => Collision_L1_n_14, A2 => Collision_L1_n_274, A3 => Collision_L1_n_315, B => Collision_L1_n_348, ZN => Collision_L1_n_367);
  Collision_L1_g14141 : NR2D0BWP7T port map(A1 => Collision_L1_n_356, A2 => Collision_L1_n_265, ZN => Collision_L1_n_366);
  Collision_L1_g14142 : OAI21D0BWP7T port map(A1 => Collision_L1_n_340, A2 => Collision_L1_n_14, B => Collision_L1_n_59, ZN => Collision_L1_n_361);
  Collision_L1_g14143 : OAI222D0BWP7T port map(A1 => Collision_L1_n_337, A2 => Collision_L1_n_302, B1 => Collision_L1_n_59, B2 => Collision_L1_n_271, C1 => Collision_L1_n_14, C2 => Collision_L1_n_270, ZN => Collision_L1_n_360);
  Collision_L1_g14144 : MAOI222D0BWP7T port map(A => Collision_L1_n_329, B => Collision_L1_n_299, C => Collision_L1_n_324, ZN => Collision_L1_n_359);
  Collision_L1_g14145 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_344, A2 => Collision_L1_n_309, B1 => Collision_L1_n_344, B2 => Collision_L1_n_309, ZN => Collision_L1_n_363);
  Collision_L1_g14146 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_326, A2 => Collision_L1_n_317, B1 => Collision_L1_n_326, B2 => Collision_L1_n_317, ZN => Collision_L1_n_362);
  Collision_L1_g14147 : OAI32D0BWP7T port map(A1 => Collision_L1_n_14, A2 => Collision_L1_n_294, A3 => Collision_L1_n_308, B1 => Collision_L1_n_293, B2 => Collision_L1_n_338, ZN => Collision_L1_n_358);
  Collision_L1_g14148 : CKND1BWP7T port map(I => Collision_L1_n_355, ZN => Collision_L1_n_356);
  Collision_L1_g14149 : CKND1BWP7T port map(I => Collision_L1_n_354, ZN => Collision_L1_n_353);
  Collision_L1_g14150 : AO21D0BWP7T port map(A1 => Collision_L1_n_333, A2 => Collision_L1_n_294, B => Collision_L1_n_342, Z => Collision_L1_n_352);
  Collision_L1_g14151 : AO211D0BWP7T port map(A1 => Collision_L1_n_274, A2 => Collision_L1_n_284, B => Collision_L1_n_331, C => Collision_L1_n_276, Z => Collision_L1_n_351);
  Collision_L1_g14152 : NR2D0BWP7T port map(A1 => Collision_L1_n_309, A2 => Collision_L1_n_341, ZN => Collision_L1_n_357);
  Collision_L1_g14153 : NR2D0BWP7T port map(A1 => Collision_L1_n_340, A2 => Collision_L1_n_263, ZN => Collision_L1_n_355);
  Collision_L1_g14154 : NR2D0BWP7T port map(A1 => Collision_L1_n_343, A2 => Collision_L1_n_287, ZN => Collision_L1_n_354);
  Collision_L1_g14155 : AOI22D0BWP7T port map(A1 => Collision_L1_n_330, A2 => Collision_L1_n_58, B1 => Collision_L1_n_280, B2 => Collision_L1_n_34, ZN => Collision_L1_n_349);
  Collision_L1_g14156 : OAI21D0BWP7T port map(A1 => Collision_L1_n_336, A2 => Collision_L1_n_34, B => Collision_L1_n_274, ZN => Collision_L1_n_348);
  Collision_L1_g14157 : OAI21D0BWP7T port map(A1 => Collision_L1_n_321, A2 => Collision_L1_n_14, B => Collision_L1_n_59, ZN => Collision_L1_n_347);
  Collision_L1_g14158 : OAI21D0BWP7T port map(A1 => Collision_L1_n_331, A2 => Collision_L1_n_14, B => Collision_L1_n_59, ZN => Collision_L1_n_346);
  Collision_L1_g14159 : IND4D0BWP7T port map(A1 => Collision_L1_n_269, B1 => Collision_L1_n_283, B2 => Collision_L1_n_316, B3 => Collision_L1_n_308, ZN => Collision_L1_n_345);
  Collision_L1_g14160 : OAI21D0BWP7T port map(A1 => Collision_L1_n_320, A2 => Collision_L1_n_286, B => Collision_L1_n_335, ZN => Collision_L1_n_350);
  Collision_L1_g14161 : HA1D0BWP7T port map(A => Collision_L1_n_3, B => Collision_L1_n_286, CO => Collision_L1_n_341, S => Collision_L1_n_344);
  Collision_L1_g14162 : ND2D0BWP7T port map(A1 => Collision_L1_n_331, A2 => Collision_L1_n_276, ZN => Collision_L1_n_343);
  Collision_L1_g14163 : NR2D0BWP7T port map(A1 => Collision_L1_n_333, A2 => Collision_L1_n_294, ZN => Collision_L1_n_342);
  Collision_L1_g14164 : IND3D0BWP7T port map(A1 => Collision_L1_n_283, B1 => Collision_L1_n_294, B2 => Collision_L1_n_314, ZN => Collision_L1_n_339);
  Collision_L1_g14165 : AOI21D0BWP7T port map(A1 => Collision_L1_n_308, A2 => Collision_L1_n_58, B => Collision_L1_n_34, ZN => Collision_L1_n_338);
  Collision_L1_g14166 : ND2D0BWP7T port map(A1 => Collision_L1_n_321, A2 => Collision_L1_n_268, ZN => Collision_L1_n_340);
  Collision_L1_g14167 : CKND1BWP7T port map(I => Collision_L1_n_335, ZN => Collision_L1_n_336);
  Collision_L1_g14168 : OR2D0BWP7T port map(A1 => Collision_L1_n_308, A2 => Collision_L1_n_314, Z => Collision_L1_n_330);
  Collision_L1_g14169 : AN2D1BWP7T port map(A1 => Collision_L1_n_307, A2 => Collision_L1_n_283, Z => Collision_L1_n_337);
  Collision_L1_g14170 : ND2D0BWP7T port map(A1 => Collision_L1_n_315, A2 => Collision_L1_n_58, ZN => Collision_L1_n_335);
  Collision_L1_g14171 : INR2D0BWP7T port map(A1 => Collision_L1_n_306, B1 => Collision_L1_n_284, ZN => Collision_L1_n_329);
  Collision_L1_g14172 : NR2D0BWP7T port map(A1 => Collision_L1_n_318, A2 => Collision_L1_n_59, ZN => Collision_L1_n_334);
  Collision_L1_g14173 : IND2D0BWP7T port map(A1 => Collision_L1_n_314, B1 => Collision_L1_n_3, ZN => Collision_L1_n_333);
  Collision_L1_g14174 : NR2D0BWP7T port map(A1 => Collision_L1_n_319, A2 => Collision_L1_n_59, ZN => Collision_L1_n_332);
  Collision_L1_g14175 : INR2D0BWP7T port map(A1 => Collision_L1_n_274, B1 => Collision_L1_n_315, ZN => Collision_L1_n_331);
  Collision_L1_g14176 : CKND1BWP7T port map(I => Collision_L1_n_323, ZN => Collision_L1_n_324);
  Collision_L1_g14177 : AOI21D0BWP7T port map(A1 => Collision_L1_n_277, A2 => Collision_L1_n_58, B => Collision_L1_n_34, ZN => Collision_L1_n_320);
  Collision_L1_g14178 : AOI21D0BWP7T port map(A1 => Collision_L1_n_277, A2 => Collision_L1_range_state_out(0), B => Collision_L1_n_309, ZN => Collision_L1_n_328);
  Collision_L1_g14179 : AOI21D0BWP7T port map(A1 => Collision_L1_n_270, A2 => Collision_L1_range_state_out(0), B => Collision_L1_n_317, ZN => Collision_L1_n_327);
  Collision_L1_g14180 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_280, A2 => Collision_L1_range_state_out(0), B1 => Collision_L1_n_280, B2 => Collision_L1_range_state_out(0), ZN => Collision_L1_n_326);
  Collision_L1_g14181 : OAI22D0BWP7T port map(A1 => Collision_L1_n_288, A2 => Collision_L1_n_3, B1 => Collision_L1_n_287, B2 => Collision_L1_range_state_out(0), ZN => Collision_L1_n_325);
  Collision_L1_g14182 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_277, A2 => Collision_L1_n_14, B1 => Collision_L1_n_277, B2 => Collision_L1_n_34, ZN => Collision_L1_n_323);
  Collision_L1_g14183 : OAI22D0BWP7T port map(A1 => Collision_L1_n_264, A2 => Collision_L1_n_3, B1 => Collision_L1_n_263, B2 => Collision_L1_range_state_out(0), ZN => Collision_L1_n_322);
  Collision_L1_g14184 : NR2D0BWP7T port map(A1 => Collision_L1_n_308, A2 => Collision_L1_n_293, ZN => Collision_L1_n_321);
  Collision_L1_g14185 : ND2D0BWP7T port map(A1 => Collision_L1_n_288, A2 => Collision_L1_n_290, ZN => Collision_L1_n_319);
  Collision_L1_g14186 : ND2D0BWP7T port map(A1 => Collision_L1_n_266, A2 => Collision_L1_n_264, ZN => Collision_L1_n_318);
  Collision_L1_g14187 : NR2D0BWP7T port map(A1 => Collision_L1_n_270, A2 => Collision_L1_range_state_out(0), ZN => Collision_L1_n_317);
  Collision_L1_g14188 : NR2D0BWP7T port map(A1 => Collision_L1_n_266, A2 => Collision_L1_n_273, ZN => Collision_L1_n_316);
  Collision_L1_g14189 : INR2D0BWP7T port map(A1 => Collision_L1_n_286, B1 => Collision_L1_n_277, ZN => Collision_L1_n_315);
  Collision_L1_g14190 : INR2D0BWP7T port map(A1 => Collision_L1_n_280, B1 => Collision_L1_n_271, ZN => Collision_L1_n_314);
  Collision_L1_g14191 : ND4D0BWP7T port map(A1 => Collision_L1_n_261, A2 => Collision_L1_n_214, A3 => Collision_L1_n_151, A4 => Collision_L1_n_110, ZN => Collision_L1_n_313);
  Collision_L1_g14192 : AN4D1BWP7T port map(A1 => Collision_L1_n_256, A2 => Collision_L1_n_215, A3 => Collision_L1_n_156, A4 => Collision_L1_n_155, Z => Collision_L1_n_312);
  Collision_L1_g14193 : AN4D1BWP7T port map(A1 => Collision_L1_n_259, A2 => Collision_L1_n_194, A3 => Collision_L1_n_139, A4 => Collision_L1_n_137, Z => Collision_L1_n_311);
  Collision_L1_g14194 : ND4D0BWP7T port map(A1 => Collision_L1_n_260, A2 => Collision_L1_n_210, A3 => Collision_L1_n_144, A4 => Collision_L1_n_123, ZN => Collision_L1_n_310);
  Collision_L1_g14195 : NR2D0BWP7T port map(A1 => Collision_L1_n_277, A2 => Collision_L1_range_state_out(0), ZN => Collision_L1_n_309);
  Collision_L1_g14196 : NR2D0BWP7T port map(A1 => Collision_L1_n_280, A2 => Collision_L1_n_270, ZN => Collision_L1_n_308);
  Collision_L1_g14197 : ND4D0BWP7T port map(A1 => Collision_L1_n_257, A2 => Collision_L1_n_204, A3 => Collision_L1_n_128, A4 => Collision_L1_n_129, ZN => Collision_L1_n_307);
  Collision_L1_g14198 : ND4D0BWP7T port map(A1 => Collision_L1_n_248, A2 => Collision_L1_n_183, A3 => Collision_L1_n_66, A4 => Collision_L1_n_67, ZN => Collision_L1_n_306);
  Collision_L1_g14199 : ND4D0BWP7T port map(A1 => Collision_L1_n_254, A2 => Collision_L1_n_197, A3 => Collision_L1_n_95, A4 => Collision_L1_n_97, ZN => Collision_L1_n_305);
  Collision_L1_g14200 : ND4D0BWP7T port map(A1 => Collision_L1_n_258, A2 => Collision_L1_n_206, A3 => Collision_L1_n_136, A4 => Collision_L1_n_131, ZN => Collision_L1_n_304);
  Collision_L1_g14201 : ND4D0BWP7T port map(A1 => Collision_L1_n_253, A2 => Collision_L1_n_195, A3 => Collision_L1_n_91, A4 => Collision_L1_n_92, ZN => Collision_L1_n_303);
  Collision_L1_g14202 : ND4D0BWP7T port map(A1 => Collision_L1_n_262, A2 => Collision_L1_n_202, A3 => Collision_L1_n_125, A4 => Collision_L1_n_126, ZN => Collision_L1_n_302);
  Collision_L1_g14203 : ND4D0BWP7T port map(A1 => Collision_L1_n_251, A2 => Collision_L1_n_191, A3 => Collision_L1_n_82, A4 => Collision_L1_n_83, ZN => Collision_L1_n_301);
  Collision_L1_g14204 : AN4D1BWP7T port map(A1 => Collision_L1_n_237, A2 => Collision_L1_n_189, A3 => Collision_L1_n_77, A4 => Collision_L1_n_78, Z => Collision_L1_n_300);
  Collision_L1_g14205 : ND4D0BWP7T port map(A1 => Collision_L1_n_249, A2 => Collision_L1_n_185, A3 => Collision_L1_n_68, A4 => Collision_L1_n_70, ZN => Collision_L1_n_299);
  Collision_L1_g14206 : ND4D0BWP7T port map(A1 => Collision_L1_n_255, A2 => Collision_L1_n_199, A3 => Collision_L1_n_105, A4 => Collision_L1_n_108, ZN => Collision_L1_n_298);
  Collision_L1_g14207 : ND4D0BWP7T port map(A1 => Collision_L1_n_247, A2 => Collision_L1_n_181, A3 => Collision_L1_n_62, A4 => Collision_L1_n_127, ZN => Collision_L1_n_297);
  Collision_L1_g14208 : AN4D1BWP7T port map(A1 => Collision_L1_n_252, A2 => Collision_L1_n_193, A3 => Collision_L1_n_86, A4 => Collision_L1_n_88, Z => Collision_L1_n_296);
  Collision_L1_g14209 : CKND1BWP7T port map(I => Collision_L1_n_294, ZN => Collision_L1_n_293);
  Collision_L1_g14210 : INVD1BWP7T port map(I => Collision_L1_n_292, ZN => Collision_L1_n_291);
  Collision_L1_g14211 : CKND1BWP7T port map(I => Collision_L1_n_290, ZN => Collision_L1_n_289);
  Collision_L1_g14212 : INVD1BWP7T port map(I => Collision_L1_n_288, ZN => Collision_L1_n_287);
  Collision_L1_g14223 : ND4D0BWP7T port map(A1 => Collision_L1_n_211, A2 => Collision_L1_n_231, A3 => Collision_L1_n_212, A4 => Collision_L1_n_119, ZN => Collision_L1_n_295);
  Collision_L1_g14224 : ND4D0BWP7T port map(A1 => Collision_L1_n_225, A2 => Collision_L1_n_118, A3 => Collision_L1_n_113, A4 => Collision_L1_n_115, ZN => Collision_L1_n_294);
  Collision_L1_g14225 : ND4D0BWP7T port map(A1 => Collision_L1_n_235, A2 => Collision_L1_n_165, A3 => Collision_L1_n_164, A4 => Collision_L1_n_167, ZN => Collision_L1_n_292);
  Collision_L1_g14226 : ND4D0BWP7T port map(A1 => Collision_L1_n_234, A2 => Collision_L1_n_160, A3 => Collision_L1_n_158, A4 => Collision_L1_n_159, ZN => Collision_L1_n_290);
  Collision_L1_g14227 : ND4D0BWP7T port map(A1 => Collision_L1_n_232, A2 => Collision_L1_n_153, A3 => Collision_L1_n_154, A4 => Collision_L1_n_152, ZN => Collision_L1_n_288);
  Collision_L1_g14228 : CKND1BWP7T port map(I => Collision_L1_n_284, ZN => Collision_L1_n_285);
  Collision_L1_g14229 : CKND1BWP7T port map(I => Collision_L1_n_281, ZN => Collision_L1_n_282);
  Collision_L1_g14231 : INVD0BWP7T port map(I => Collision_L1_n_276, ZN => Collision_L1_n_275);
  Collision_L1_g14232 : CKND1BWP7T port map(I => Collision_L1_n_273, ZN => Collision_L1_n_272);
  Collision_L1_g14233 : CKND1BWP7T port map(I => Collision_L1_n_270, ZN => Collision_L1_n_271);
  Collision_L1_g14234 : INVD0BWP7T port map(I => Collision_L1_n_268, ZN => Collision_L1_n_267);
  Collision_L1_g14235 : INVD1BWP7T port map(I => Collision_L1_n_266, ZN => Collision_L1_n_265);
  Collision_L1_g14236 : INVD1BWP7T port map(I => Collision_L1_n_264, ZN => Collision_L1_n_263);
  Collision_L1_g14237 : AN4D1BWP7T port map(A1 => Collision_L1_n_228, A2 => Collision_L1_n_134, A3 => Collision_L1_n_121, A4 => Collision_L1_n_133, Z => Collision_L1_n_286);
  Collision_L1_g14238 : ND4D0BWP7T port map(A1 => Collision_L1_n_226, A2 => Collision_L1_n_116, A3 => Collision_L1_n_117, A4 => Collision_L1_n_114, ZN => Collision_L1_n_284);
  Collision_L1_g14239 : AN4D1BWP7T port map(A1 => Collision_L1_n_221, A2 => Collision_L1_n_87, A3 => Collision_L1_n_84, A4 => Collision_L1_n_85, Z => Collision_L1_n_283);
  Collision_L1_g14240 : ND4D0BWP7T port map(A1 => Collision_L1_n_187, A2 => Collision_L1_n_219, A3 => Collision_L1_n_186, A4 => Collision_L1_n_145, ZN => Collision_L1_n_281);
  Collision_L1_g14241 : ND4D0BWP7T port map(A1 => Collision_L1_n_224, A2 => Collision_L1_n_107, A3 => Collision_L1_n_109, A4 => Collision_L1_n_106, ZN => Collision_L1_n_280);
  Collision_L1_g14242 : ND4D0BWP7T port map(A1 => Collision_L1_n_217, A2 => Collision_L1_n_64, A3 => Collision_L1_n_65, A4 => Collision_L1_n_63, ZN => Collision_L1_n_278);
  Collision_L1_g14243 : ND4D0BWP7T port map(A1 => Collision_L1_n_227, A2 => Collision_L1_n_122, A3 => Collision_L1_n_146, A4 => Collision_L1_n_161, ZN => Collision_L1_n_277);
  Collision_L1_g14244 : ND4D0BWP7T port map(A1 => Collision_L1_n_230, A2 => Collision_L1_n_179, A3 => Collision_L1_n_147, A4 => Collision_L1_n_149, ZN => Collision_L1_n_276);
  Collision_L1_g14245 : ND4D0BWP7T port map(A1 => Collision_L1_n_229, A2 => Collision_L1_n_141, A3 => Collision_L1_n_142, A4 => Collision_L1_n_138, ZN => Collision_L1_n_274);
  Collision_L1_g14246 : ND4D0BWP7T port map(A1 => Collision_L1_n_220, A2 => Collision_L1_n_79, A3 => Collision_L1_n_76, A4 => Collision_L1_n_80, ZN => Collision_L1_n_273);
  Collision_L1_g14247 : ND4D0BWP7T port map(A1 => Collision_L1_n_223, A2 => Collision_L1_n_101, A3 => Collision_L1_n_103, A4 => Collision_L1_n_100, ZN => Collision_L1_n_270);
  Collision_L1_g14248 : ND4D0BWP7T port map(A1 => Collision_L1_n_222, A2 => Collision_L1_n_94, A3 => Collision_L1_n_96, A4 => Collision_L1_n_93, ZN => Collision_L1_n_269);
  Collision_L1_g14249 : ND4D0BWP7T port map(A1 => Collision_L1_n_209, A2 => Collision_L1_n_102, A3 => Collision_L1_n_162, A4 => Collision_L1_n_140, ZN => Collision_L1_n_268);
  Collision_L1_g14250 : ND4D0BWP7T port map(A1 => Collision_L1_n_218, A2 => Collision_L1_n_74, A3 => Collision_L1_n_71, A4 => Collision_L1_n_73, ZN => Collision_L1_n_266);
  Collision_L1_g14251 : ND4D0BWP7T port map(A1 => Collision_L1_n_233, A2 => Collision_L1_n_124, A3 => Collision_L1_n_132, A4 => Collision_L1_n_166, ZN => Collision_L1_n_264);
  Collision_L1_g14252 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => x_pos_e2(1), B1 => Collision_L1_n_32, B2 => x_pos_e1(1), C => Collision_L1_n_201, ZN => Collision_L1_n_262);
  Collision_L1_g14253 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => x_pos_e2(4), B1 => Collision_L1_n_32, B2 => x_pos_e1(4), C => Collision_L1_n_213, ZN => Collision_L1_n_261);
  Collision_L1_g14254 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => x_pos_e2(6), B1 => Collision_L1_n_32, B2 => x_pos_e1(6), C => Collision_L1_n_236, ZN => Collision_L1_n_260);
  Collision_L1_g14255 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => x_pos_e2(3), B1 => Collision_L1_n_32, B2 => x_pos_e1(3), C => Collision_L1_n_207, ZN => Collision_L1_n_259);
  Collision_L1_g14256 : AOI221D0BWP7T port map(A1 => Collision_L1_n_49, A2 => x_pos_b3(2), B1 => Collision_L1_n_4, B2 => x_pos_p(2), C => Collision_L1_n_205, ZN => Collision_L1_n_258);
  Collision_L1_g14257 : AOI221D0BWP7T port map(A1 => Collision_L1_n_46, A2 => x_pos_e6(0), B1 => Collision_L1_n_47, B2 => x_pos_e5(0), C => Collision_L1_n_203, ZN => Collision_L1_n_257);
  Collision_L1_g14258 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => x_pos_e2(7), B1 => Collision_L1_n_32, B2 => x_pos_e1(7), C => Collision_L1_n_200, ZN => Collision_L1_n_256);
  Collision_L1_g14259 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => y_pos_e2(8), B1 => Collision_L1_n_32, B2 => y_pos_e1(8), C => Collision_L1_n_198, ZN => Collision_L1_n_255);
  Collision_L1_g14260 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => y_pos_e2(4), B1 => Collision_L1_n_32, B2 => y_pos_e1(4), C => Collision_L1_n_196, ZN => Collision_L1_n_254);
  Collision_L1_g14261 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => y_pos_e2(5), B1 => Collision_L1_n_32, B2 => y_pos_e1(5), C => Collision_L1_n_208, ZN => Collision_L1_n_253);
  Collision_L1_g14262 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => y_pos_e2(7), B1 => Collision_L1_n_32, B2 => y_pos_e1(7), C => Collision_L1_n_192, ZN => Collision_L1_n_252);
  Collision_L1_g14263 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => y_pos_e2(6), B1 => Collision_L1_n_32, B2 => y_pos_e1(6), C => Collision_L1_n_190, ZN => Collision_L1_n_251);
  Collision_L1_g14265 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_56, A2 => Collision_L1_n_30, B1 => Collision_L1_n_169, B2 => collision_output_vector(14), ZN => Collision_L1_n_250);
  Collision_L1_g14266 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => y_pos_e2(1), B1 => Collision_L1_n_32, B2 => y_pos_e1(1), C => Collision_L1_n_184, ZN => Collision_L1_n_249);
  Collision_L1_g14267 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => y_pos_e2(0), B1 => Collision_L1_n_32, B2 => y_pos_e1(0), C => Collision_L1_n_182, ZN => Collision_L1_n_248);
  Collision_L1_g14268 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => x_pos_e2(8), B1 => Collision_L1_n_32, B2 => x_pos_e1(8), C => Collision_L1_n_180, ZN => Collision_L1_n_247);
  Collision_L1_g14269 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_56, A2 => Collision_L1_n_6, B1 => Collision_L1_n_177, B2 => collision_output_vector(4), ZN => Collision_L1_n_246);
  Collision_L1_g14270 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_56, A2 => Collision_L1_n_28, B1 => Collision_L1_n_178, B2 => collision_output_vector(1), ZN => Collision_L1_n_245);
  Collision_L1_g14271 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_56, A2 => Collision_L1_n_41, B1 => Collision_L1_n_176, B2 => collision_output_vector(10), ZN => Collision_L1_n_244);
  Collision_L1_g14272 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_56, A2 => Collision_L1_n_45, B1 => Collision_L1_n_175, B2 => collision_output_vector(11), ZN => Collision_L1_n_243);
  Collision_L1_g14273 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_56, A2 => Collision_L1_n_18, B1 => Collision_L1_n_174, B2 => collision_output_vector(12), ZN => Collision_L1_n_242);
  Collision_L1_g14274 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_56, A2 => Collision_L1_n_39, B1 => Collision_L1_n_173, B2 => collision_output_vector(13), ZN => Collision_L1_n_241);
  Collision_L1_g14275 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_56, A2 => Collision_L1_n_36, B1 => Collision_L1_n_172, B2 => collision_output_vector(2), ZN => Collision_L1_n_240);
  Collision_L1_g14276 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_56, A2 => Collision_L1_n_42, B1 => Collision_L1_n_171, B2 => collision_output_vector(9), ZN => Collision_L1_n_239);
  Collision_L1_g14277 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_56, A2 => Collision_L1_n_15, B1 => Collision_L1_n_170, B2 => collision_output_vector(0), ZN => Collision_L1_n_238);
  Collision_L1_g14278 : AOI221D0BWP7T port map(A1 => Collision_L1_n_33, A2 => y_pos_e2(3), B1 => Collision_L1_n_32, B2 => y_pos_e1(3), C => Collision_L1_n_188, ZN => Collision_L1_n_237);
  Collision_L1_g14279 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => x_pos_e4(6), B1 => x_pos_e3(6), B2 => Collision_L1_n_51, Z => Collision_L1_n_236);
  Collision_L1_g14280 : AOI221D0BWP7T port map(A1 => Collision_L1_n_29, A2 => y_pos_b2(7), B1 => Collision_L1_n_16, B2 => y_pos_b1(7), C => Collision_L1_n_163, ZN => Collision_L1_n_235);
  Collision_L1_g14281 : AOI221D0BWP7T port map(A1 => Collision_L1_n_44, A2 => y_pos_e3(6), B1 => Collision_L1_n_17, B2 => y_pos_e4(6), C => Collision_L1_n_157, ZN => Collision_L1_n_234);
  Collision_L1_g14282 : AOI221D0BWP7T port map(A1 => Collision_L1_n_29, A2 => x_pos_b2(5), B1 => Collision_L1_n_16, B2 => x_pos_b1(5), C => Collision_L1_n_89, ZN => Collision_L1_n_233);
  Collision_L1_g14283 : AOI221D0BWP7T port map(A1 => Collision_L1_n_29, A2 => y_pos_b2(5), B1 => Collision_L1_n_16, B2 => y_pos_b1(5), C => Collision_L1_n_150, ZN => Collision_L1_n_232);
  Collision_L1_g14284 : AOI221D0BWP7T port map(A1 => Collision_L1_n_46, A2 => x_pos_e6(5), B1 => Collision_L1_n_4, B2 => x_pos_p(5), C => Collision_L1_n_148, ZN => Collision_L1_n_231);
  Collision_L1_g14285 : AOI221D0BWP7T port map(A1 => Collision_L1_n_29, A2 => y_pos_b2(4), B1 => Collision_L1_n_16, B2 => y_pos_b1(4), C => Collision_L1_n_143, ZN => Collision_L1_n_230);
  Collision_L1_g14286 : AOI221D0BWP7T port map(A1 => Collision_L1_n_29, A2 => y_pos_b2(3), B1 => Collision_L1_n_16, B2 => y_pos_b1(3), C => Collision_L1_n_135, ZN => Collision_L1_n_229);
  Collision_L1_g14287 : AOI221D0BWP7T port map(A1 => Collision_L1_n_44, A2 => y_pos_e3(2), B1 => Collision_L1_n_17, B2 => y_pos_e4(2), C => Collision_L1_n_130, ZN => Collision_L1_n_228);
  Collision_L1_g14288 : AOI221D0BWP7T port map(A1 => Collision_L1_n_29, A2 => y_pos_b2(1), B1 => Collision_L1_n_16, B2 => y_pos_b1(1), C => Collision_L1_n_98, ZN => Collision_L1_n_227);
  Collision_L1_g14289 : AOI221D0BWP7T port map(A1 => Collision_L1_n_29, A2 => y_pos_b2(0), B1 => Collision_L1_n_16, B2 => y_pos_b1(0), C => Collision_L1_n_112, ZN => Collision_L1_n_226);
  Collision_L1_g14290 : AOI221D0BWP7T port map(A1 => Collision_L1_n_44, A2 => x_pos_e3(3), B1 => Collision_L1_n_17, B2 => x_pos_e4(3), C => Collision_L1_n_111, ZN => Collision_L1_n_225);
  Collision_L1_g14291 : AOI221D0BWP7T port map(A1 => Collision_L1_n_29, A2 => x_pos_b2(2), B1 => Collision_L1_n_16, B2 => x_pos_b1(2), C => Collision_L1_n_104, ZN => Collision_L1_n_224);
  Collision_L1_g14292 : AOI221D0BWP7T port map(A1 => Collision_L1_n_29, A2 => x_pos_b2(1), B1 => Collision_L1_n_16, B2 => x_pos_b1(1), C => Collision_L1_n_99, ZN => Collision_L1_n_223);
  Collision_L1_g14293 : AOI221D0BWP7T port map(A1 => Collision_L1_n_44, A2 => x_pos_e3(8), B1 => Collision_L1_n_17, B2 => x_pos_e4(8), C => Collision_L1_n_120, ZN => Collision_L1_n_222);
  Collision_L1_g14294 : AOI221D0BWP7T port map(A1 => Collision_L1_n_44, A2 => x_pos_e3(0), B1 => Collision_L1_n_17, B2 => x_pos_e4(0), C => Collision_L1_n_81, ZN => Collision_L1_n_221);
  Collision_L1_g14295 : AOI221D0BWP7T port map(A1 => Collision_L1_n_29, A2 => x_pos_b2(7), B1 => Collision_L1_n_16, B2 => x_pos_b1(7), C => Collision_L1_n_75, ZN => Collision_L1_n_220);
  Collision_L1_g14296 : AOI221D0BWP7T port map(A1 => Collision_L1_n_46, A2 => y_pos_e6(2), B1 => Collision_L1_n_4, B2 => y_pos_p(2), C => Collision_L1_n_72, ZN => Collision_L1_n_219);
  Collision_L1_g14297 : AOI221D0BWP7T port map(A1 => Collision_L1_n_44, A2 => x_pos_e3(6), B1 => Collision_L1_n_17, B2 => x_pos_e4(6), C => Collision_L1_n_69, ZN => Collision_L1_n_218);
  Collision_L1_g14298 : AOI221D0BWP7T port map(A1 => Collision_L1_n_29, A2 => y_pos_b2(8), B1 => Collision_L1_n_16, B2 => y_pos_b1(8), C => Collision_L1_n_61, ZN => Collision_L1_n_217);
  Collision_L1_g14299 : OAI22D0BWP7T port map(A1 => Collision_L1_n_15, A2 => Collision_L1_n_50, B1 => Collision_L1_n_55, B2 => reset, ZN => Collision_L1_n_216);
  Collision_L1_g14300 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => x_pos_b1(7), B1 => Collision_L1_n_48, B2 => x_pos_b2(7), ZN => Collision_L1_n_215);
  Collision_L1_g14301 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => x_pos_b1(4), B1 => Collision_L1_n_48, B2 => x_pos_b2(4), ZN => Collision_L1_n_214);
  Collision_L1_g14302 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => x_pos_e4(4), B1 => x_pos_e3(4), B2 => Collision_L1_n_51, Z => Collision_L1_n_213);
  Collision_L1_g14303 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => x_pos_b1(5), B1 => Collision_L1_n_48, B2 => x_pos_b2(5), ZN => Collision_L1_n_212);
  Collision_L1_g14304 : AOI22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => x_pos_e4(5), B1 => Collision_L1_n_51, B2 => x_pos_e3(5), ZN => Collision_L1_n_211);
  Collision_L1_g14305 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => x_pos_b1(6), B1 => Collision_L1_n_48, B2 => x_pos_b2(6), ZN => Collision_L1_n_210);
  Collision_L1_g14306 : AOI221D0BWP7T port map(A1 => Collision_L1_n_44, A2 => x_pos_e3(4), B1 => Collision_L1_n_17, B2 => x_pos_e4(4), C => Collision_L1_n_90, ZN => Collision_L1_n_209);
  Collision_L1_g14307 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => y_pos_e4(5), B1 => y_pos_e3(5), B2 => Collision_L1_n_51, Z => Collision_L1_n_208);
  Collision_L1_g14308 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => x_pos_e4(3), B1 => x_pos_e3(3), B2 => Collision_L1_n_51, Z => Collision_L1_n_207);
  Collision_L1_g14309 : AOI22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => x_pos_e4(2), B1 => Collision_L1_n_51, B2 => x_pos_e3(2), ZN => Collision_L1_n_206);
  Collision_L1_g14310 : AO22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => x_pos_b1(2), B1 => x_pos_b2(2), B2 => Collision_L1_n_48, Z => Collision_L1_n_205);
  Collision_L1_g14311 : AOI22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => x_pos_e4(0), B1 => Collision_L1_n_51, B2 => x_pos_e3(0), ZN => Collision_L1_n_204);
  Collision_L1_g14312 : AO22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => x_pos_b1(0), B1 => x_pos_b2(0), B2 => Collision_L1_n_48, Z => Collision_L1_n_203);
  Collision_L1_g14313 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => x_pos_b1(1), B1 => Collision_L1_n_48, B2 => x_pos_b2(1), ZN => Collision_L1_n_202);
  Collision_L1_g14314 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => x_pos_e4(1), B1 => x_pos_e3(1), B2 => Collision_L1_n_51, Z => Collision_L1_n_201);
  Collision_L1_g14315 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => x_pos_e4(7), B1 => x_pos_e3(7), B2 => Collision_L1_n_51, Z => Collision_L1_n_200);
  Collision_L1_g14316 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => y_pos_b1(8), B1 => Collision_L1_n_48, B2 => y_pos_b2(8), ZN => Collision_L1_n_199);
  Collision_L1_g14317 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => y_pos_e4(8), B1 => y_pos_e3(8), B2 => Collision_L1_n_51, Z => Collision_L1_n_198);
  Collision_L1_g14318 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => y_pos_b1(4), B1 => Collision_L1_n_48, B2 => y_pos_b2(4), ZN => Collision_L1_n_197);
  Collision_L1_g14319 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => y_pos_e4(4), B1 => y_pos_e3(4), B2 => Collision_L1_n_51, Z => Collision_L1_n_196);
  Collision_L1_g14320 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => y_pos_b1(5), B1 => Collision_L1_n_48, B2 => y_pos_b2(5), ZN => Collision_L1_n_195);
  Collision_L1_g14321 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => x_pos_b1(3), B1 => Collision_L1_n_48, B2 => x_pos_b2(3), ZN => Collision_L1_n_194);
  Collision_L1_g14322 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => y_pos_b1(7), B1 => Collision_L1_n_48, B2 => y_pos_b2(7), ZN => Collision_L1_n_193);
  Collision_L1_g14323 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => y_pos_e4(7), B1 => y_pos_e3(7), B2 => Collision_L1_n_51, Z => Collision_L1_n_192);
  Collision_L1_g14324 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => y_pos_b1(6), B1 => Collision_L1_n_48, B2 => y_pos_b2(6), ZN => Collision_L1_n_191);
  Collision_L1_g14325 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => y_pos_e4(6), B1 => y_pos_e3(6), B2 => Collision_L1_n_51, Z => Collision_L1_n_190);
  Collision_L1_g14326 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => y_pos_b1(3), B1 => Collision_L1_n_48, B2 => y_pos_b2(3), ZN => Collision_L1_n_189);
  Collision_L1_g14327 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => y_pos_e4(3), B1 => y_pos_e3(3), B2 => Collision_L1_n_51, Z => Collision_L1_n_188);
  Collision_L1_g14328 : AOI22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => y_pos_e4(2), B1 => Collision_L1_n_51, B2 => y_pos_e3(2), ZN => Collision_L1_n_187);
  Collision_L1_g14329 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => y_pos_b1(2), B1 => Collision_L1_n_48, B2 => y_pos_b2(2), ZN => Collision_L1_n_186);
  Collision_L1_g14330 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => y_pos_b1(1), B1 => Collision_L1_n_48, B2 => y_pos_b2(1), ZN => Collision_L1_n_185);
  Collision_L1_g14331 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => y_pos_e4(1), B1 => y_pos_e3(1), B2 => Collision_L1_n_51, Z => Collision_L1_n_184);
  Collision_L1_g14332 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => y_pos_b1(0), B1 => Collision_L1_n_48, B2 => y_pos_b2(0), ZN => Collision_L1_n_183);
  Collision_L1_g14333 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => y_pos_e4(0), B1 => y_pos_e3(0), B2 => Collision_L1_n_51, Z => Collision_L1_n_182);
  Collision_L1_g14334 : AOI22D0BWP7T port map(A1 => Collision_L1_n_52, A2 => x_pos_b1(8), B1 => Collision_L1_n_48, B2 => x_pos_b2(8), ZN => Collision_L1_n_181);
  Collision_L1_g14335 : AO22D0BWP7T port map(A1 => Collision_L1_n_53, A2 => x_pos_e4(8), B1 => x_pos_e3(8), B2 => Collision_L1_n_51, Z => Collision_L1_n_180);
  Collision_L1_g14336 : AOI22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => y_pos_e2(4), B1 => Collision_L1_n_43, B2 => y_pos_e1(4), ZN => Collision_L1_n_179);
  Collision_L1_g14337 : OAI21D0BWP7T port map(A1 => Collision_L1_n_29, A2 => reset, B => Collision_L1_n_57, ZN => Collision_L1_n_178);
  Collision_L1_g14338 : OAI21D0BWP7T port map(A1 => Collision_L1_n_484, A2 => reset, B => Collision_L1_n_57, ZN => Collision_L1_n_177);
  Collision_L1_g14339 : OAI21D0BWP7T port map(A1 => Collision_L1_n_40, A2 => reset, B => Collision_L1_n_57, ZN => Collision_L1_n_176);
  Collision_L1_g14340 : OAI21D0BWP7T port map(A1 => Collision_L1_n_44, A2 => reset, B => Collision_L1_n_57, ZN => Collision_L1_n_175);
  Collision_L1_g14341 : OAI21D0BWP7T port map(A1 => Collision_L1_n_17, A2 => reset, B => Collision_L1_n_57, ZN => Collision_L1_n_174);
  Collision_L1_g14342 : OAI21D0BWP7T port map(A1 => Collision_L1_n_38, A2 => reset, B => Collision_L1_n_57, ZN => Collision_L1_n_173);
  Collision_L1_g14343 : OAI21D0BWP7T port map(A1 => Collision_L1_n_37, A2 => reset, B => Collision_L1_n_57, ZN => Collision_L1_n_172);
  Collision_L1_g14344 : OAI21D0BWP7T port map(A1 => Collision_L1_n_43, A2 => reset, B => Collision_L1_n_57, ZN => Collision_L1_n_171);
  Collision_L1_g14345 : OAI21D0BWP7T port map(A1 => Collision_L1_n_16, A2 => reset, B => Collision_L1_n_57, ZN => Collision_L1_n_170);
  Collision_L1_g14346 : OAI21D0BWP7T port map(A1 => Collision_L1_n_31, A2 => reset, B => Collision_L1_n_57, ZN => Collision_L1_n_169);
  Collision_L1_g14347 : OAI32D0BWP7T port map(A1 => Collision_L1_n_5, A2 => Collision_L1_n_7, A3 => Collision_L1_n_8, B1 => Collision_L1_n_9, B2 => Collision_start_value_s(0), ZN => Collision_L1_n_168);
  Collision_L1_g14348 : AOI22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => y_pos_e5(7), B1 => Collision_L1_n_31, B2 => y_pos_e6(7), ZN => Collision_L1_n_167);
  Collision_L1_g14349 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => x_pos_b3(5), B1 => Collision_L1_n_484, B2 => x_pos_p(5), ZN => Collision_L1_n_166);
  Collision_L1_g14350 : AOI22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => y_pos_e2(7), B1 => Collision_L1_n_43, B2 => y_pos_e1(7), ZN => Collision_L1_n_165);
  Collision_L1_g14351 : AOI22D0BWP7T port map(A1 => Collision_L1_n_44, A2 => y_pos_e3(7), B1 => Collision_L1_n_17, B2 => y_pos_e4(7), ZN => Collision_L1_n_164);
  Collision_L1_g14352 : AO22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => y_pos_b3(7), B1 => y_pos_p(7), B2 => Collision_L1_n_484, Z => Collision_L1_n_163);
  Collision_L1_g14353 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => x_pos_b3(4), B1 => Collision_L1_n_484, B2 => x_pos_p(4), ZN => Collision_L1_n_162);
  Collision_L1_g14354 : AOI22D0BWP7T port map(A1 => Collision_L1_n_44, A2 => y_pos_e3(1), B1 => Collision_L1_n_17, B2 => y_pos_e4(1), ZN => Collision_L1_n_161);
  Collision_L1_g14355 : AOI22D0BWP7T port map(A1 => Collision_L1_n_29, A2 => y_pos_b2(6), B1 => Collision_L1_n_16, B2 => y_pos_b1(6), ZN => Collision_L1_n_160);
  Collision_L1_g14356 : AOI22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => y_pos_e5(6), B1 => Collision_L1_n_31, B2 => y_pos_e6(6), ZN => Collision_L1_n_159);
  Collision_L1_g14357 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => y_pos_b3(6), B1 => Collision_L1_n_484, B2 => y_pos_p(6), ZN => Collision_L1_n_158);
  Collision_L1_g14358 : AO22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => y_pos_e2(6), B1 => y_pos_e1(6), B2 => Collision_L1_n_43, Z => Collision_L1_n_157);
  Collision_L1_g14359 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => x_pos_e6(7), B1 => Collision_L1_n_47, B2 => x_pos_e5(7), ZN => Collision_L1_n_156);
  Collision_L1_g14360 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => x_pos_b3(7), B1 => Collision_L1_n_4, B2 => x_pos_p(7), ZN => Collision_L1_n_155);
  Collision_L1_g14361 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => y_pos_b3(5), B1 => Collision_L1_n_484, B2 => y_pos_p(5), ZN => Collision_L1_n_154);
  Collision_L1_g14362 : AOI22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => y_pos_e2(5), B1 => Collision_L1_n_43, B2 => y_pos_e1(5), ZN => Collision_L1_n_153);
  Collision_L1_g14363 : AOI22D0BWP7T port map(A1 => Collision_L1_n_44, A2 => y_pos_e3(5), B1 => Collision_L1_n_17, B2 => y_pos_e4(5), ZN => Collision_L1_n_152);
  Collision_L1_g14364 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => x_pos_b3(4), B1 => Collision_L1_n_47, B2 => x_pos_e5(4), ZN => Collision_L1_n_151);
  Collision_L1_g14365 : AO22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => y_pos_e5(5), B1 => y_pos_e6(5), B2 => Collision_L1_n_31, Z => Collision_L1_n_150);
  Collision_L1_g14366 : AOI22D0BWP7T port map(A1 => Collision_L1_n_44, A2 => y_pos_e3(4), B1 => Collision_L1_n_17, B2 => y_pos_e4(4), ZN => Collision_L1_n_149);
  Collision_L1_g14367 : AO22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => x_pos_b3(5), B1 => x_pos_e5(5), B2 => Collision_L1_n_47, Z => Collision_L1_n_148);
  Collision_L1_g14368 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => y_pos_b3(4), B1 => Collision_L1_n_484, B2 => y_pos_p(4), ZN => Collision_L1_n_147);
  Collision_L1_g14369 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => y_pos_b3(1), B1 => Collision_L1_n_484, B2 => y_pos_p(1), ZN => Collision_L1_n_146);
  Collision_L1_g14370 : AOI22D0BWP7T port map(A1 => Collision_L1_n_33, A2 => y_pos_e2(2), B1 => Collision_L1_n_32, B2 => y_pos_e1(2), ZN => Collision_L1_n_145);
  Collision_L1_g14371 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => x_pos_e6(6), B1 => Collision_L1_n_47, B2 => x_pos_e5(6), ZN => Collision_L1_n_144);
  Collision_L1_g14372 : AO22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => y_pos_e5(4), B1 => y_pos_e6(4), B2 => Collision_L1_n_31, Z => Collision_L1_n_143);
  Collision_L1_g14373 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => y_pos_b3(3), B1 => Collision_L1_n_484, B2 => y_pos_p(3), ZN => Collision_L1_n_142);
  Collision_L1_g14374 : AOI22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => y_pos_e2(3), B1 => Collision_L1_n_43, B2 => y_pos_e1(3), ZN => Collision_L1_n_141);
  Collision_L1_g14375 : AOI22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => x_pos_e5(4), B1 => Collision_L1_n_31, B2 => x_pos_e6(4), ZN => Collision_L1_n_140);
  Collision_L1_g14376 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => x_pos_e6(3), B1 => Collision_L1_n_47, B2 => x_pos_e5(3), ZN => Collision_L1_n_139);
  Collision_L1_g14377 : AOI22D0BWP7T port map(A1 => Collision_L1_n_44, A2 => y_pos_e3(3), B1 => Collision_L1_n_17, B2 => y_pos_e4(3), ZN => Collision_L1_n_138);
  Collision_L1_g14378 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => x_pos_b3(3), B1 => Collision_L1_n_4, B2 => x_pos_p(3), ZN => Collision_L1_n_137);
  Collision_L1_g14379 : AOI22D0BWP7T port map(A1 => Collision_L1_n_33, A2 => x_pos_e2(2), B1 => Collision_L1_n_32, B2 => x_pos_e1(2), ZN => Collision_L1_n_136);
  Collision_L1_g14380 : AO22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => y_pos_e5(3), B1 => y_pos_e6(3), B2 => Collision_L1_n_31, Z => Collision_L1_n_135);
  Collision_L1_g14381 : AOI22D0BWP7T port map(A1 => Collision_L1_n_29, A2 => y_pos_b2(2), B1 => Collision_L1_n_16, B2 => y_pos_b1(2), ZN => Collision_L1_n_134);
  Collision_L1_g14382 : AOI22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => y_pos_e5(2), B1 => Collision_L1_n_31, B2 => y_pos_e6(2), ZN => Collision_L1_n_133);
  Collision_L1_g14383 : AOI22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => x_pos_e2(5), B1 => Collision_L1_n_43, B2 => x_pos_e1(5), ZN => Collision_L1_n_132);
  Collision_L1_g14384 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => x_pos_e6(2), B1 => Collision_L1_n_47, B2 => x_pos_e5(2), ZN => Collision_L1_n_131);
  Collision_L1_g14385 : AO22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => y_pos_e2(2), B1 => y_pos_e1(2), B2 => Collision_L1_n_43, Z => Collision_L1_n_130);
  Collision_L1_g14386 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => x_pos_b3(0), B1 => Collision_L1_n_4, B2 => x_pos_p(0), ZN => Collision_L1_n_129);
  Collision_L1_g14387 : AOI22D0BWP7T port map(A1 => Collision_L1_n_33, A2 => x_pos_e2(0), B1 => Collision_L1_n_32, B2 => x_pos_e1(0), ZN => Collision_L1_n_128);
  Collision_L1_g14388 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => x_pos_e6(8), B1 => Collision_L1_n_4, B2 => x_pos_p(8), ZN => Collision_L1_n_127);
  Collision_L1_g14389 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => x_pos_e6(1), B1 => Collision_L1_n_4, B2 => x_pos_p(1), ZN => Collision_L1_n_126);
  Collision_L1_g14390 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => x_pos_b3(1), B1 => Collision_L1_n_47, B2 => x_pos_e5(1), ZN => Collision_L1_n_125);
  Collision_L1_g14391 : AOI22D0BWP7T port map(A1 => Collision_L1_n_44, A2 => x_pos_e3(5), B1 => Collision_L1_n_17, B2 => x_pos_e4(5), ZN => Collision_L1_n_124);
  Collision_L1_g14392 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => x_pos_b3(6), B1 => Collision_L1_n_4, B2 => x_pos_p(6), ZN => Collision_L1_n_123);
  Collision_L1_g14393 : AOI22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => y_pos_e2(1), B1 => Collision_L1_n_43, B2 => y_pos_e1(1), ZN => Collision_L1_n_122);
  Collision_L1_g14394 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => y_pos_b3(2), B1 => Collision_L1_n_484, B2 => y_pos_p(2), ZN => Collision_L1_n_121);
  Collision_L1_g14396 : AO22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => x_pos_e2(8), B1 => x_pos_e1(8), B2 => Collision_L1_n_43, Z => Collision_L1_n_120);
  Collision_L1_g14397 : AOI22D0BWP7T port map(A1 => Collision_L1_n_33, A2 => x_pos_e2(5), B1 => Collision_L1_n_32, B2 => x_pos_e1(5), ZN => Collision_L1_n_119);
  Collision_L1_g14398 : AOI22D0BWP7T port map(A1 => Collision_L1_n_29, A2 => x_pos_b2(3), B1 => Collision_L1_n_16, B2 => x_pos_b1(3), ZN => Collision_L1_n_118);
  Collision_L1_g14399 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => y_pos_b3(0), B1 => Collision_L1_n_484, B2 => y_pos_p(0), ZN => Collision_L1_n_117);
  Collision_L1_g14400 : AOI22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => y_pos_e2(0), B1 => Collision_L1_n_43, B2 => y_pos_e1(0), ZN => Collision_L1_n_116);
  Collision_L1_g14401 : AOI22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => x_pos_e5(3), B1 => Collision_L1_n_31, B2 => x_pos_e6(3), ZN => Collision_L1_n_115);
  Collision_L1_g14402 : AOI22D0BWP7T port map(A1 => Collision_L1_n_44, A2 => y_pos_e3(0), B1 => Collision_L1_n_17, B2 => y_pos_e4(0), ZN => Collision_L1_n_114);
  Collision_L1_g14403 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => x_pos_b3(3), B1 => Collision_L1_n_484, B2 => x_pos_p(3), ZN => Collision_L1_n_113);
  Collision_L1_g14404 : AO22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => y_pos_e5(0), B1 => y_pos_e6(0), B2 => Collision_L1_n_31, Z => Collision_L1_n_112);
  Collision_L1_g14405 : AO22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => x_pos_e2(3), B1 => x_pos_e1(3), B2 => Collision_L1_n_43, Z => Collision_L1_n_111);
  Collision_L1_g14406 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => x_pos_e6(4), B1 => Collision_L1_n_4, B2 => x_pos_p(4), ZN => Collision_L1_n_110);
  Collision_L1_g14407 : AOI22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => x_pos_e2(2), B1 => Collision_L1_n_43, B2 => x_pos_e1(2), ZN => Collision_L1_n_109);
  Collision_L1_g14408 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => y_pos_b3(8), B1 => Collision_L1_n_4, B2 => y_pos_p(8), ZN => Collision_L1_n_108);
  Collision_L1_g14409 : AOI22D0BWP7T port map(A1 => Collision_L1_n_44, A2 => x_pos_e3(2), B1 => Collision_L1_n_17, B2 => x_pos_e4(2), ZN => Collision_L1_n_107);
  Collision_L1_g14410 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => x_pos_b3(2), B1 => Collision_L1_n_484, B2 => x_pos_p(2), ZN => Collision_L1_n_106);
  Collision_L1_g14411 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => y_pos_e6(8), B1 => Collision_L1_n_47, B2 => y_pos_e5(8), ZN => Collision_L1_n_105);
  Collision_L1_g14412 : AO22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => x_pos_e5(2), B1 => x_pos_e6(2), B2 => Collision_L1_n_31, Z => Collision_L1_n_104);
  Collision_L1_g14413 : AOI22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => x_pos_e2(1), B1 => Collision_L1_n_43, B2 => x_pos_e1(1), ZN => Collision_L1_n_103);
  Collision_L1_g14414 : AOI22D0BWP7T port map(A1 => Collision_L1_n_29, A2 => x_pos_b2(4), B1 => Collision_L1_n_16, B2 => x_pos_b1(4), ZN => Collision_L1_n_102);
  Collision_L1_g14415 : AOI22D0BWP7T port map(A1 => Collision_L1_n_44, A2 => x_pos_e3(1), B1 => Collision_L1_n_17, B2 => x_pos_e4(1), ZN => Collision_L1_n_101);
  Collision_L1_g14416 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => x_pos_b3(1), B1 => Collision_L1_n_484, B2 => x_pos_p(1), ZN => Collision_L1_n_100);
  Collision_L1_g14417 : AO22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => x_pos_e5(1), B1 => x_pos_e6(1), B2 => Collision_L1_n_31, Z => Collision_L1_n_99);
  Collision_L1_g14418 : AO22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => y_pos_e5(1), B1 => y_pos_e6(1), B2 => Collision_L1_n_31, Z => Collision_L1_n_98);
  Collision_L1_g14419 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => y_pos_b3(4), B1 => Collision_L1_n_4, B2 => y_pos_p(4), ZN => Collision_L1_n_97);
  Collision_L1_g14420 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => x_pos_b3(8), B1 => Collision_L1_n_484, B2 => x_pos_p(8), ZN => Collision_L1_n_96);
  Collision_L1_g14421 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => y_pos_e6(4), B1 => Collision_L1_n_47, B2 => y_pos_e5(4), ZN => Collision_L1_n_95);
  Collision_L1_g14422 : AOI22D0BWP7T port map(A1 => Collision_L1_n_29, A2 => x_pos_b2(8), B1 => Collision_L1_n_16, B2 => x_pos_b1(8), ZN => Collision_L1_n_94);
  Collision_L1_g14423 : AOI22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => x_pos_e5(8), B1 => Collision_L1_n_31, B2 => x_pos_e6(8), ZN => Collision_L1_n_93);
  Collision_L1_g14424 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => y_pos_e6(5), B1 => Collision_L1_n_4, B2 => y_pos_p(5), ZN => Collision_L1_n_92);
  Collision_L1_g14425 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => y_pos_b3(5), B1 => Collision_L1_n_47, B2 => y_pos_e5(5), ZN => Collision_L1_n_91);
  Collision_L1_g14426 : AO22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => x_pos_e2(4), B1 => x_pos_e1(4), B2 => Collision_L1_n_43, Z => Collision_L1_n_90);
  Collision_L1_g14427 : AO22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => x_pos_e5(5), B1 => x_pos_e6(5), B2 => Collision_L1_n_31, Z => Collision_L1_n_89);
  Collision_L1_g14428 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => y_pos_b3(7), B1 => Collision_L1_n_4, B2 => y_pos_p(7), ZN => Collision_L1_n_88);
  Collision_L1_g14429 : AOI22D0BWP7T port map(A1 => Collision_L1_n_29, A2 => x_pos_b2(0), B1 => Collision_L1_n_16, B2 => x_pos_b1(0), ZN => Collision_L1_n_87);
  Collision_L1_g14430 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => y_pos_e6(7), B1 => Collision_L1_n_47, B2 => y_pos_e5(7), ZN => Collision_L1_n_86);
  Collision_L1_g14431 : AOI22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => x_pos_e5(0), B1 => Collision_L1_n_31, B2 => x_pos_e6(0), ZN => Collision_L1_n_85);
  Collision_L1_g14432 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => x_pos_b3(0), B1 => Collision_L1_n_484, B2 => x_pos_p(0), ZN => Collision_L1_n_84);
  Collision_L1_g14433 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => y_pos_e6(6), B1 => Collision_L1_n_4, B2 => y_pos_p(6), ZN => Collision_L1_n_83);
  Collision_L1_g14434 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => y_pos_b3(6), B1 => Collision_L1_n_47, B2 => y_pos_e5(6), ZN => Collision_L1_n_82);
  Collision_L1_g14435 : AO22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => x_pos_e2(0), B1 => x_pos_e1(0), B2 => Collision_L1_n_43, Z => Collision_L1_n_81);
  Collision_L1_g14436 : AOI22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => x_pos_e5(7), B1 => Collision_L1_n_31, B2 => x_pos_e6(7), ZN => Collision_L1_n_80);
  Collision_L1_g14437 : AOI22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => x_pos_e2(7), B1 => Collision_L1_n_43, B2 => x_pos_e1(7), ZN => Collision_L1_n_79);
  Collision_L1_g14438 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => y_pos_e6(3), B1 => Collision_L1_n_4, B2 => y_pos_p(3), ZN => Collision_L1_n_78);
  Collision_L1_g14439 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => y_pos_b3(3), B1 => Collision_L1_n_47, B2 => y_pos_e5(3), ZN => Collision_L1_n_77);
  Collision_L1_g14440 : AOI22D0BWP7T port map(A1 => Collision_L1_n_44, A2 => x_pos_e3(7), B1 => Collision_L1_n_17, B2 => x_pos_e4(7), ZN => Collision_L1_n_76);
  Collision_L1_g14441 : AO22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => x_pos_b3(7), B1 => x_pos_p(7), B2 => Collision_L1_n_484, Z => Collision_L1_n_75);
  Collision_L1_g14442 : AOI22D0BWP7T port map(A1 => Collision_L1_n_29, A2 => x_pos_b2(6), B1 => Collision_L1_n_16, B2 => x_pos_b1(6), ZN => Collision_L1_n_74);
  Collision_L1_g14443 : AOI22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => x_pos_e5(6), B1 => Collision_L1_n_31, B2 => x_pos_e6(6), ZN => Collision_L1_n_73);
  Collision_L1_g14444 : AO22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => y_pos_b3(2), B1 => y_pos_e5(2), B2 => Collision_L1_n_47, Z => Collision_L1_n_72);
  Collision_L1_g14445 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => x_pos_b3(6), B1 => Collision_L1_n_484, B2 => x_pos_p(6), ZN => Collision_L1_n_71);
  Collision_L1_g14446 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => y_pos_b3(1), B1 => Collision_L1_n_4, B2 => y_pos_p(1), ZN => Collision_L1_n_70);
  Collision_L1_g14447 : AO22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => x_pos_e2(6), B1 => x_pos_e1(6), B2 => Collision_L1_n_43, Z => Collision_L1_n_69);
  Collision_L1_g14448 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => y_pos_e6(1), B1 => Collision_L1_n_47, B2 => y_pos_e5(1), ZN => Collision_L1_n_68);
  Collision_L1_g14449 : AOI22D0BWP7T port map(A1 => Collision_L1_n_46, A2 => y_pos_e6(0), B1 => Collision_L1_n_4, B2 => y_pos_p(0), ZN => Collision_L1_n_67);
  Collision_L1_g14450 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => y_pos_b3(0), B1 => Collision_L1_n_47, B2 => y_pos_e5(0), ZN => Collision_L1_n_66);
  Collision_L1_g14451 : AOI22D0BWP7T port map(A1 => Collision_L1_n_40, A2 => y_pos_e2(8), B1 => Collision_L1_n_43, B2 => y_pos_e1(8), ZN => Collision_L1_n_65);
  Collision_L1_g14452 : AOI22D0BWP7T port map(A1 => Collision_L1_n_44, A2 => y_pos_e3(8), B1 => Collision_L1_n_17, B2 => y_pos_e4(8), ZN => Collision_L1_n_64);
  Collision_L1_g14453 : AOI22D0BWP7T port map(A1 => Collision_L1_n_37, A2 => y_pos_b3(8), B1 => Collision_L1_n_484, B2 => y_pos_p(8), ZN => Collision_L1_n_63);
  Collision_L1_g14454 : AOI22D0BWP7T port map(A1 => Collision_L1_n_49, A2 => x_pos_b3(8), B1 => Collision_L1_n_47, B2 => x_pos_e5(8), ZN => Collision_L1_n_62);
  Collision_L1_g14455 : AO22D0BWP7T port map(A1 => Collision_L1_n_38, A2 => y_pos_e5(8), B1 => y_pos_e6(8), B2 => Collision_L1_n_31, Z => Collision_L1_n_61);
  Collision_L1_g14456 : ND4D0BWP7T port map(A1 => Collision_L1_n_25, A2 => Collision_L1_n_26, A3 => Collision_L1_n_27, A4 => Collision_L1_n_23, ZN => Collision_L1_n_60);
  Collision_L1_g14457 : INVD1BWP7T port map(I => Collision_L1_n_34, ZN => Collision_L1_n_59);
  Collision_L1_g14458 : INVD1BWP7T port map(I => Collision_L1_n_14, ZN => Collision_L1_n_58);
  Collision_L1_g14459 : IND2D0BWP7T port map(A1 => Collision_L1_n_35, B1 => Collision_L1_state(2), ZN => Collision_L1_n_55);
  Collision_L1_g14460 : ND2D0BWP7T port map(A1 => Collision_L1_n_50, A2 => Collision_L1_n_1, ZN => Collision_L1_n_57);
  Collision_L1_g14461 : OR2D0BWP7T port map(A1 => Collision_L1_n_50, A2 => Collision_L1_state(0), Z => Collision_L1_n_56);
  Collision_L1_g14462 : IND3D0BWP7T port map(A1 => Collision_enable_s, B1 => Collision_L1_state(0), B2 => Collision_L1_n_22, ZN => Collision_L1_n_54);
  Collision_L1_g14463 : NR3D0BWP7T port map(A1 => Collision_L1_n_8, A2 => Collision_count_2_s(0), A3 => Collision_count_2_s(1), ZN => Collision_L1_n_53);
  Collision_L1_g14464 : AN3D0BWP7T port map(A1 => Collision_L1_n_9, A2 => Collision_L1_n_7, A3 => Collision_L1_n_5, Z => Collision_L1_n_52);
  Collision_L1_g14465 : NR3D0BWP7T port map(A1 => Collision_L1_n_10, A2 => Collision_L1_n_7, A3 => Collision_L1_n_5, ZN => Collision_L1_n_51);
  Collision_L1_g14466 : INVD1BWP7T port map(I => Collision_L1_n_44, ZN => Collision_L1_n_45);
  Collision_L1_g14467 : INVD1BWP7T port map(I => Collision_L1_n_43, ZN => Collision_L1_n_42);
  Collision_L1_g14468 : INVD1BWP7T port map(I => Collision_L1_n_40, ZN => Collision_L1_n_41);
  Collision_L1_g14469 : INVD1BWP7T port map(I => Collision_L1_n_38, ZN => Collision_L1_n_39);
  Collision_L1_g14470 : INVD1BWP7T port map(I => Collision_L1_n_37, ZN => Collision_L1_n_36);
  Collision_L1_g14471 : ND2D0BWP7T port map(A1 => Collision_L1_n_22, A2 => Collision_enable_s, ZN => Collision_L1_n_50);
  Collision_L1_g14472 : INR2D0BWP7T port map(A1 => Collision_L1_n_9, B1 => Collision_L1_n_19, ZN => Collision_L1_n_49);
  Collision_L1_g14473 : INR2D0BWP7T port map(A1 => Collision_L1_n_9, B1 => Collision_L1_n_13, ZN => Collision_L1_n_48);
  Collision_L1_g14474 : NR2D0BWP7T port map(A1 => Collision_L1_n_8, A2 => Collision_L1_n_13, ZN => Collision_L1_n_47);
  Collision_L1_g14475 : NR2D0BWP7T port map(A1 => Collision_L1_n_19, A2 => Collision_L1_n_8, ZN => Collision_L1_n_46);
  Collision_L1_g14476 : NR2D0BWP7T port map(A1 => Collision_L1_n_20, A2 => Collision_L1_n_11, ZN => Collision_L1_n_44);
  Collision_L1_g14477 : NR2D0BWP7T port map(A1 => Collision_L1_n_501, A2 => Collision_L1_n_11, ZN => Collision_L1_n_43);
  Collision_L1_g14478 : NR2D0BWP7T port map(A1 => Collision_L1_n_503, A2 => Collision_L1_n_20, ZN => Collision_L1_n_40);
  Collision_L1_g14479 : NR2D0BWP7T port map(A1 => Collision_L1_n_502, A2 => Collision_L1_n_11, ZN => Collision_L1_n_38);
  Collision_L1_g14480 : NR2D0BWP7T port map(A1 => Collision_L1_n_500, A2 => Collision_L1_n_20, ZN => Collision_L1_n_37);
  Collision_L1_g14481 : INVD1BWP7T port map(I => Collision_L1_n_30, ZN => Collision_L1_n_31);
  Collision_L1_g14482 : INVD1BWP7T port map(I => Collision_L1_n_29, ZN => Collision_L1_n_28);
  Collision_L1_g14483 : XNR2D1BWP7T port map(A1 => Collision_count_2_s(3), A2 => Collision_count_1_s(3), ZN => Collision_L1_n_27);
  Collision_L1_g14484 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_5, A2 => Collision_count_1_s(0), B1 => Collision_L1_n_5, B2 => Collision_count_1_s(0), ZN => Collision_L1_n_26);
  Collision_L1_g14485 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_7, A2 => Collision_count_1_s(1), B1 => Collision_L1_n_7, B2 => Collision_count_1_s(1), ZN => Collision_L1_n_25);
  Collision_L1_g14486 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_483, A2 => Collision_L1_n_482, B1 => Collision_L1_n_6, B2 => Collision_L1_n_481, ZN => Collision_L1_n_24);
  Collision_L1_g14487 : XNR2D1BWP7T port map(A1 => Collision_count_2_s(2), A2 => Collision_count_1_s(2), ZN => Collision_L1_n_23);
  Collision_L1_g14488 : IND3D0BWP7T port map(A1 => Collision_enable_s, B1 => n_5, B2 => Collision_L1_n_2, ZN => Collision_L1_n_35);
  Collision_L1_g14489 : MOAI22D0BWP7T port map(A1 => Collision_L1_n_3, A2 => Collision_L1_range_state_out(1), B1 => Collision_L1_n_3, B2 => Collision_L1_range_state_out(1), ZN => Collision_L1_n_34);
  Collision_L1_g14490 : NR2D0BWP7T port map(A1 => Collision_L1_n_19, A2 => Collision_L1_n_10, ZN => Collision_L1_n_33);
  Collision_L1_g14491 : NR2D0BWP7T port map(A1 => Collision_L1_n_13, A2 => Collision_L1_n_10, ZN => Collision_L1_n_32);
  Collision_L1_g14492 : IND3D0BWP7T port map(A1 => Collision_L1_n_503, B1 => Collision_count_1_s(1), B2 => Collision_count_1_s(2), ZN => Collision_L1_n_30);
  Collision_L1_g14493 : INR3D0BWP7T port map(A1 => Collision_count_1_s(0), B1 => Collision_count_1_s(3), B2 => Collision_L1_n_501, ZN => Collision_L1_n_29);
  Collision_L1_g14494 : CKND1BWP7T port map(I => Collision_L1_n_22, ZN => Collision_L1_n_21);
  Collision_L1_g14495 : INVD1BWP7T port map(I => Collision_L1_n_17, ZN => Collision_L1_n_18);
  Collision_L1_g14496 : INVD1BWP7T port map(I => Collision_L1_n_16, ZN => Collision_L1_n_15);
  Collision_L1_g14497 : NR2D0BWP7T port map(A1 => Collision_L1_state(2), A2 => reset, ZN => Collision_L1_n_22);
  Collision_L1_g14498 : IND2D0BWP7T port map(A1 => Collision_count_1_s(2), B1 => Collision_count_1_s(1), ZN => Collision_L1_n_20);
  Collision_L1_g14499 : ND2D0BWP7T port map(A1 => Collision_L1_n_5, A2 => Collision_count_2_s(1), ZN => Collision_L1_n_19);
  Collision_L1_g14500 : NR2D0BWP7T port map(A1 => Collision_L1_n_503, A2 => Collision_L1_n_502, ZN => Collision_L1_n_17);
  Collision_L1_g14501 : NR2D0BWP7T port map(A1 => Collision_L1_n_500, A2 => Collision_L1_n_501, ZN => Collision_L1_n_16);
  Collision_L1_g14502 : ND2D0BWP7T port map(A1 => Collision_L1_range_state_out(0), A2 => Collision_L1_range_state_out(1), ZN => Collision_L1_n_14);
  Collision_L1_g14503 : ND2D0BWP7T port map(A1 => Collision_L1_n_7, A2 => Collision_count_2_s(0), ZN => Collision_L1_n_13);
  Collision_L1_g14504 : IND2D0BWP7T port map(A1 => Collision_L1_range_state_out(1), B1 => Collision_L1_n_3, ZN => Collision_L1_n_12);
  Collision_L1_g14505 : ND2D0BWP7T port map(A1 => Collision_count_1_s(0), A2 => Collision_count_1_s(3), ZN => Collision_L1_n_11);
  Collision_L1_g14506 : IND2D0BWP7T port map(A1 => Collision_count_2_s(2), B1 => Collision_count_2_s(3), ZN => Collision_L1_n_10);
  Collision_L1_g14507 : NR2D0BWP7T port map(A1 => Collision_count_2_s(2), A2 => Collision_count_2_s(3), ZN => Collision_L1_n_9);
  Collision_L1_g14508 : ND2D0BWP7T port map(A1 => Collision_count_2_s(3), A2 => Collision_count_2_s(2), ZN => Collision_L1_n_8);
  Collision_L1_g14509 : INVD1BWP7T port map(I => Collision_count_2_s(1), ZN => Collision_L1_n_7);
  Collision_L1_g14511 : INVD1BWP7T port map(I => Collision_L1_n_484, ZN => Collision_L1_n_6);
  Collision_L1_g14513 : INVD1BWP7T port map(I => Collision_count_2_s(0), ZN => Collision_L1_n_5);
  Collision_L1_range_state_out_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => Collision_L1_n_1, D => Collision_L1_n_24, Q => Collision_L1_range_state_out(0), QN => Collision_L1_n_3);
  Collision_L1_drc_bufs14517 : INVD0BWP7T port map(I => reset, ZN => Collision_L1_n_1);
  Collision_L1_g2 : NR2D1BWP7T port map(A1 => Collision_L1_n_504, A2 => Collision_L1_n_269, ZN => Collision_L1_n_505);
  Collision_L1_g3 : OA21D0BWP7T port map(A1 => Collision_L1_n_334, A2 => Collision_L1_n_366, B => Collision_L1_n_273, Z => Collision_L1_n_504);
  Collision_L1_g14524 : IND3D1BWP7T port map(A1 => Collision_L1_n_278, B1 => Collision_L1_n_509, B2 => Collision_L1_n_12, ZN => Collision_L1_n_506);
  Collision_L1_g14526 : IOA22D0BWP7T port map(A1 => Collision_L1_n_476, A2 => Collision_count_1_s(2), B1 => Collision_L1_n_501, B2 => Collision_L1_n_503, ZN => Collision_start_value_s(2));
  Collision_L1_g14527 : MAOI22D0BWP7T port map(A1 => Collision_L1_n_332, A2 => Collision_L1_n_292, B1 => Collision_L1_n_369, B2 => Collision_L1_n_291, ZN => Collision_L1_n_509);
  Collision_L2_count_inside_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => Collision_L2_n_1, D => Collision_L2_n_8, Q => Collision_count_1_s(3));
  Collision_L2_count_inside_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => Collision_L2_n_1, D => Collision_L2_n_7, Q => Collision_count_1_s(2));
  Collision_L2_g71 : MOAI22D0BWP7T port map(A1 => Collision_L2_n_6, A2 => Collision_count_1_s(3), B1 => Collision_L2_n_6, B2 => Collision_count_1_s(3), ZN => Collision_L2_n_8);
  Collision_L2_count_inside_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => Collision_L2_n_1, D => Collision_L2_n_5, Q => Collision_count_1_s(1));
  Collision_L2_g73 : MOAI22D0BWP7T port map(A1 => Collision_L2_n_4, A2 => Collision_count_1_s(2), B1 => Collision_L2_n_4, B2 => Collision_count_1_s(2), ZN => Collision_L2_n_7);
  Collision_L2_g74 : IND2D0BWP7T port map(A1 => Collision_L2_n_4, B1 => Collision_count_1_s(2), ZN => Collision_L2_n_6);
  Collision_L2_count_inside_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => Collision_L2_n_1, D => Collision_L2_n_3, Q => Collision_count_1_s(0));
  Collision_L2_g76 : MOAI22D0BWP7T port map(A1 => Collision_L2_n_2, A2 => Collision_count_1_s(1), B1 => Collision_L2_n_2, B2 => Collision_count_1_s(1), ZN => Collision_L2_n_5);
  Collision_L2_g77 : IND2D0BWP7T port map(A1 => Collision_L2_n_2, B1 => Collision_count_1_s(1), ZN => Collision_L2_n_4);
  Collision_L2_g78 : CKXOR2D0BWP7T port map(A1 => Collision_count_1_s(0), A2 => Collision_enable_s, Z => Collision_L2_n_3);
  Collision_L2_g79 : ND2D0BWP7T port map(A1 => Collision_enable_s, A2 => Collision_count_1_s(0), ZN => Collision_L2_n_2);
  Collision_L2_g80 : INVD1BWP7T port map(I => reset, ZN => Collision_L2_n_1);
  Collision_L3_count_inside_reg_3 : DFND1BWP7T port map(CPN => clk, D => Collision_L3_n_13, Q => Collision_count_2_s(3), QN => UNCONNECTED3);
  Collision_L3_g182 : AO22D0BWP7T port map(A1 => Collision_L3_n_11, A2 => Collision_L3_n_5, B1 => Collision_start_value_s(3), B2 => Collision_L3_n_3, Z => Collision_L3_n_13);
  Collision_L3_count_inside_reg_2 : DFND1BWP7T port map(CPN => clk, D => Collision_L3_n_12, Q => Collision_count_2_s(2), QN => UNCONNECTED4);
  Collision_L3_g184 : AO22D0BWP7T port map(A1 => Collision_L3_n_10, A2 => Collision_L3_n_5, B1 => Collision_L3_n_3, B2 => Collision_start_value_s(2), Z => Collision_L3_n_12);
  Collision_L3_g185 : MOAI22D0BWP7T port map(A1 => Collision_L3_n_9, A2 => Collision_count_2_s(3), B1 => Collision_L3_n_9, B2 => Collision_count_2_s(3), ZN => Collision_L3_n_11);
  Collision_L3_count_inside_reg_1 : DFND1BWP7T port map(CPN => clk, D => Collision_L3_n_8, Q => Collision_count_2_s(1), QN => UNCONNECTED5);
  Collision_L3_g187 : MOAI22D0BWP7T port map(A1 => Collision_L3_n_4, A2 => Collision_count_2_s(2), B1 => Collision_L3_n_4, B2 => Collision_count_2_s(2), ZN => Collision_L3_n_10);
  Collision_L3_count_inside_reg_0 : DFND1BWP7T port map(CPN => clk, D => Collision_L3_n_7, Q => Collision_count_2_s(0), QN => Collision_L3_n_2);
  Collision_L3_g189 : INR2D0BWP7T port map(A1 => Collision_L3_n_5, B1 => Collision_L3_n_6, ZN => Collision_L3_n_8);
  Collision_L3_g190 : IND2D0BWP7T port map(A1 => Collision_L3_n_4, B1 => Collision_count_2_s(2), ZN => Collision_L3_n_9);
  Collision_L3_g191 : AO22D0BWP7T port map(A1 => Collision_L3_n_5, A2 => Collision_L3_n_2, B1 => Collision_L3_n_3, B2 => Collision_start_value_s(0), Z => Collision_L3_n_7);
  Collision_L3_g192 : MAOI22D0BWP7T port map(A1 => Collision_L3_n_2, A2 => Collision_count_2_s(1), B1 => Collision_L3_n_2, B2 => Collision_count_2_s(1), ZN => Collision_L3_n_6);
  Collision_L3_g193 : NR2D0BWP7T port map(A1 => Collision_reset_2_s, A2 => reset, ZN => Collision_L3_n_5);
  Collision_L3_g194 : ND2D0BWP7T port map(A1 => Collision_count_2_s(0), A2 => Collision_count_2_s(1), ZN => Collision_L3_n_4);
  Collision_L3_g195 : INR2D0BWP7T port map(A1 => Collision_reset_2_s, B1 => reset, ZN => Collision_L3_n_3);

end synthesised;
