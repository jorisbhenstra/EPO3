library IEEE;
use IEEE.std_logic_1164.ALL;

entity col_top_level_tb is
end col_top_level_tb;

