configuration spawn_timer_behaviour_cfg of spawn_timer is
   for behaviour
   end for;
end spawn_timer_behaviour_cfg;
