configuration state_gradius_behaviour_cfg of state_gradius is
   for behaviour
   end for;
end state_gradius_behaviour_cfg;
